* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XANTENNA__8507__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7257__I1 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7963_ _0189_ net156 mod.Data_Mem.F_M.MRAM\[779\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5968__A1 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7009__I1 mod.Data_Mem.F_M.MRAM\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6914_ _3253_ mod.Data_Mem.F_M.MRAM\[13\]\[5\] _3381_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7894_ _0120_ net205 mod.Data_Mem.F_M.MRAM\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4640__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6845_ _3256_ mod.Data_Mem.F_M.MRAM\[769\]\[6\] _3340_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6776_ _3297_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3988_ mod.Arithmetic.ACTI.x\[0\] _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8499__D _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8515_ _0019_ net355 mod.Data_Mem.F_M.out_data\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5727_ mod.Data_Mem.F_M.MRAM\[14\]\[0\] mod.Data_Mem.F_M.MRAM\[15\]\[0\] _2351_ _2352_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7256__I _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8446_ _0542_ net373 mod.Data_Mem.F_M.MRAM\[793\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6145__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5658_ _2054_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4609_ _1159_ _1196_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8377_ _0473_ net316 mod.Data_Mem.F_M.MRAM\[784\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _2224_ mod.Data_Mem.F_M.MRAM\[31\]\[4\] mod.Data_Mem.F_M.MRAM\[30\]\[4\] _2225_
+ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7328_ _3297_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8126__RN net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6448__A2 mod.Data_Mem.F_M.MRAM\[780\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7259_ mod.Data_Mem.F_M.MRAM\[31\]\[5\] _3316_ _3590_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4459__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8187__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7248__I1 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3959__I _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4056__S _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4631__A1 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6384__A1 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5187__A2 mod.Data_Mem.F_M.MRAM\[771\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6136__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7487__I1 mod.Data_Mem.F_M.MRAM\[781\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5414__I _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6298__S1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout260_I net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout358_I net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _1539_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4622__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4891_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _3205_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6375__A1 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6561_ mod.Data_Mem.F_M.MRAM\[781\]\[7\] _3115_ _3005_ mod.Data_Mem.F_M.MRAM\[769\]\[7\]
+ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7076__I mod.Data_Mem.F_M.MRAM\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8300_ _0396_ net95 mod.Data_Mem.F_M.MRAM\[773\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5512_ _1547_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6127__A1 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ mod.Data_Mem.F_M.MRAM\[12\]\[4\] mod.Data_Mem.F_M.MRAM\[14\]\[4\] mod.Data_Mem.F_M.MRAM\[13\]\[4\]
+ _1870_ _2273_ _2500_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8231_ mod.P1.instr_reg\[17\] net23 net240 mod.P2.dest_reg1\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5443_ _1727_ _2091_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4689__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8162_ mod.Data_Mem.F_M.out_data\[72\] net30 net270 mod.Arithmetic.I_out\[72\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5374_ mod.Data_Mem.F_M.MRAM\[771\]\[7\] mod.Data_Mem.F_M.MRAM\[770\]\[7\] _1906_
+ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5350__A2 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7113_ _3504_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8108__RN net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7478__I1 mod.Data_Mem.F_M.MRAM\[780\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4325_ _0994_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout105 net108 net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_8093_ mod.Data_Mem.F_M.out_data\[3\] net56 net336 mod.Arithmetic.ACTI.x\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout116 net117 net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout127 net129 net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout138 net141 net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _3468_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout149 net151 net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ _0828_ _0930_ _0660_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4187_ _0629_ _0855_ _0862_ mod.P3.Res\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6989__I0 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7946_ _0172_ net88 mod.Data_Mem.F_M.MRAM\[789\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7877_ _0103_ net376 mod.Data_Mem.F_M.MRAM\[24\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6828_ mod.Data_Mem.F_M.dest\[1\] _3333_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6366__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _3286_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__I1 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6118__A1 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7166__I0 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8429_ _0525_ net162 mod.Data_Mem.F_M.MRAM\[791\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4144__A3 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5234__I _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__S _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__I _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__I3 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5409__I _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7157__I0 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout106_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__I1 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ mod.Arithmetic.ACTI.x\[4\] _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ _1500_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4041_ _0690_ _0717_ _0708_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5891__I0 mod.Data_Mem.F_M.MRAM\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7800_ _3898_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5992_ _2136_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5399__A2 _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7731_ _3859_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4943_ mod.Data_Mem.F_M.MRAM\[787\]\[0\] mod.Data_Mem.F_M.MRAM\[786\]\[0\] _1611_
+ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4071__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6703__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7662_ mod.Data_Mem.F_M.MRAM\[790\]\[7\] _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4874_ _1542_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6613_ mod.Data_Mem.F_M.MRAM\[24\]\[2\] _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7593_ _3786_ _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_fanout19_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5020__A1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4223__I mod.Arithmetic.CN.I_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6544_ _3145_ _3146_ _2425_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7148__I0 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _3002_ _3080_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8214_ _0315_ net150 mod.Data_Mem.F_M.MRAM\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5426_ _2080_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6520__A1 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8145_ mod.Data_Mem.F_M.out_data\[55\] net63 net361 mod.Arithmetic.CN.I_in\[55\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5357_ mod.Data_Mem.F_M.MRAM\[15\]\[7\] _1886_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7470__S _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4098__C _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _0980_ _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_82_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8076_ mod.P3.Res\[4\] net34 net261 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__7320__I0 _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5288_ mod.Data_Mem.F_M.MRAM\[773\]\[5\] mod.Data_Mem.F_M.MRAM\[772\]\[5\] _1876_
+ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7027_ _3447_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4239_ _0846_ _0912_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_56_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__B1 _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8225__CLK net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7929_ _0155_ net368 mod.Data_Mem.F_M.MRAM\[8\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4062__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6339__A1 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8375__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7139__I0 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3972__I _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5078__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6578__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5139__I _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout223_I net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _1039_ _1144_ _1147_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5553__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6260_ _1661_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6502__A1 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5305__A2 mod.Data_Mem.F_M.MRAM\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _1873_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__7892__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6191_ _2744_ _2802_ _2805_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _1644_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5069__A1 mod.Data_Mem.F_M.MRAM\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5073_ _1575_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4024_ mod.Arithmetic.CN.I_in\[22\] _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4292__A2 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__I1 mod.Data_Mem.F_M.MRAM\[786\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5975_ _2351_ _1938_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7714_ mod.Data_Mem.F_M.MRAM\[794\]\[1\] _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4926_ _1594_ _1552_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7645_ _3816_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4857_ _1525_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5049__I _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7576_ _3749_ mod.Data_Mem.F_M.MRAM\[785\]\[2\] _3773_ _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5544__A2 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _1235_ _1344_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6527_ _3049_ _3130_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4888__I _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ _2057_ _3064_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4355__I0 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5409_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6389_ _2247_ _2250_ _2995_ _2998_ _1489_ _2784_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_88_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8128_ mod.Data_Mem.F_M.out_data\[38\] net44 net251 mod.Arithmetic.CN.I_in\[38\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8059_ _0268_ net95 mod.Data_Mem.F_M.MRAM\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5512__I _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4283__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3967__I _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A2 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6032__I0 mod.Data_Mem.F_M.MRAM\[770\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5535__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7780__I0 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5299__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout173_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4038__I mod.Arithmetic.CN.I_in\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5074__I1 mod.Data_Mem.F_M.MRAM\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7763__A3 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout340_I net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _2203_ _2380_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4711_ _1369_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _2289_ mod.Data_Mem.F_M.MRAM\[29\]\[5\] _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7285__S _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7430_ _3688_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4642_ _1311_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7771__I0 _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7361_ mod.Data_Mem.F_M.MRAM\[772\]\[5\] _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4573_ _0640_ mod.Arithmetic.ACTI.x\[5\] _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7084__I mod.Data_Mem.F_M.MRAM\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6312_ _1657_ _1953_ _2870_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7292_ _3305_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6487__B1 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6243_ _2854_ _2214_ _2855_ _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6487__C2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8070__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6174_ _2209_ mod.Data_Mem.F_M.MRAM\[783\]\[2\] mod.Data_Mem.F_M.MRAM\[782\]\[2\]
+ _2280_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5125_ _1518_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ _1508_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4007_ mod.Arithmetic.CN.I_in\[21\] _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5958_ _2570_ _2576_ _2577_ _2258_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4909_ mod.Data_Mem.F_M.MRAM\[774\]\[0\] _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5889_ mod.Data_Mem.F_M.MRAM\[4\]\[3\] mod.Data_Mem.F_M.MRAM\[5\]\[3\] mod.Data_Mem.F_M.MRAM\[20\]\[3\]
+ mod.Data_Mem.F_M.MRAM\[21\]\[3\] _1796_ _1757_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7628_ _3319_ _3798_ _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5935__C _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7559_ _3765_ mod.Data_Mem.F_M.MRAM\[784\]\[3\] _3760_ _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8563__CLK net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4059__S _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_404 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_415 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_426 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_437 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_448 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_459 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A1 _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4256__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__A2 mod.Data_Mem.F_M.MRAM\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8093__CLK net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4192__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7505__I0 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7632__I mod.Data_Mem.F_M.MRAM\[788\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout290_I net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout388_I net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5819__I0 mod.Data_Mem.F_M.MRAM\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7930__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5444__A1 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__I0 mod.Data_Mem.F_M.MRAM\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5295__I1 mod.Data_Mem.F_M.MRAM\[770\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6930_ _3394_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5995__A2 mod.Data_Mem.F_M.MRAM\[773\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6861_ mod.Data_Mem.F_M.MRAM\[779\]\[6\] _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7197__A1 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8115__D mod.Data_Mem.F_M.out_data\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5812_ _2432_ _2433_ _2435_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6792_ _3310_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8531_ _0035_ net328 mod.Data_Mem.F_M.out_data\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5743_ _1594_ _1501_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6711__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8462_ _0558_ net384 mod.Data_Mem.F_M.MRAM\[795\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5674_ _1904_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7413_ mod.Data_Mem.F_M.MRAM\[775\]\[7\] _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4625_ _1292_ _0743_ _1295_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8393_ _0489_ net201 mod.Data_Mem.F_M.MRAM\[786\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7344_ _3315_ _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4556_ _0643_ mod.Arithmetic.CN.I_in\[58\] mod.Arithmetic.CN.I_in\[59\] _1136_ _1228_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__8586__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7275_ mod.Data_Mem.F_M.MRAM\[5\]\[5\] _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4487_ _1089_ _1102_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _2827_ _2830_ _2831_ _2091_ _2839_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6158__I _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ _1558_ _1705_ _1707_ _2772_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5108_ mod.Data_Mem.F_M.MRAM\[768\]\[2\] _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ _1873_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ mod.Data_Mem.F_M.MRAM\[775\]\[1\] mod.Data_Mem.F_M.MRAM\[774\]\[1\] _1706_
+ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A2 mod.Data_Mem.F_M.MRAM\[788\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3997__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__B _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5237__I mod.Data_Mem.F_M.MRAM\[783\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4141__I _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4174__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5910__A2 mod.Data_Mem.F_M.MRAM\[786\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput7 net7 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__B1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_fanout136_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5147__I _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7563__S _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout303_I net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4051__I mod.Arithmetic.CN.I_in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4410_ _1048_ _1077_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4165__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5390_ _2033_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4704__A3 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4341_ _1008_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ mod.Data_Mem.F_M.MRAM\[20\]\[1\] _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout309 net310 net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4272_ _0869_ _0887_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6701__I1 mod.Data_Mem.F_M.MRAM\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5665__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4468__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6011_ _2548_ _2623_ _2626_ _2629_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7962_ _0188_ net316 mod.Data_Mem.F_M.MRAM\[779\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5968__A2 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6090__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6913_ _3382_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout49_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7893_ _0119_ net383 mod.Data_Mem.F_M.MRAM\[25\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6217__I0 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4640__A2 mod.Arithmetic.CN.I_in\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6844_ _1955_ _3337_ _3344_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4670__B _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6775_ mod.Data_Mem.F_M.dest\[8\] mod.DMen_reg2 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3987_ _0661_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8071__RN net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6441__I _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8514_ _0018_ net331 mod.Data_Mem.F_M.out_data\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5726_ _1695_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8445_ _0541_ net377 mod.Data_Mem.F_M.MRAM\[793\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5657_ _2164_ _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7473__S _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4156__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _1162_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7976__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5588_ _1815_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8376_ _0472_ net215 mod.Data_Mem.F_M.MRAM\[784\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4896__I _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7327_ _3633_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4539_ mod.Arithmetic.CN.I_in\[43\] _1096_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7258_ _3591_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6209_ _2820_ _2821_ _2822_ _2823_ _2679_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7189_ _3523_ mod.Data_Mem.F_M.MRAM\[29\]\[0\] _3550_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4631__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4395__A1 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4698__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5647__A1 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__I1 mod.Data_Mem.F_M.MRAM\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8281__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout253_I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4890_ _1534_ _1558_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4386__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7999__CLK net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _2827_ _3161_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5511_ _2118_ _2150_ _2152_ _2132_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6491_ _2345_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5806__S _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4138__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8230_ mod.P1.instr_reg\[13\] net17 net223 mod.P2.dest_reg1\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5442_ _2090_ _1622_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5886__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4689__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5373_ mod.Data_Mem.F_M.MRAM\[769\]\[7\] mod.Data_Mem.F_M.MRAM\[768\]\[7\] _1904_
+ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8161_ mod.Data_Mem.F_M.out_data\[71\] net62 net358 mod.Arithmetic.CN.I_in\[71\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__7092__I mod.Data_Mem.F_M.MRAM\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7112_ _3452_ mod.Data_Mem.F_M.MRAM\[3\]\[2\] _3501_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4324_ _0930_ _0995_ _0996_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8092_ mod.Data_Mem.F_M.out_data\[2\] net59 net348 mod.Arithmetic.ACTI.x\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout106 net108 net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout117 net120 net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5638__A1 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7043_ _3450_ mod.Data_Mem.F_M.MRAM\[1\]\[1\] _3466_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout128 net129 net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout139 net141 net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4255_ mod.Arithmetic.CN.I_in\[49\] _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4186_ _0754_ _0857_ _0859_ _0861_ _0628_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6989__I1 mod.Data_Mem.F_M.MRAM\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7945_ _0171_ net142 mod.Data_Mem.F_M.MRAM\[789\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7468__S _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7876_ _0102_ net386 mod.Data_Mem.F_M.MRAM\[24\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6827_ mod.Data_Mem.F_M.dest\[0\] _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6366__A2 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8004__CLK net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6758_ mod.Data_Mem.F_M.MRAM\[8\]\[2\] _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5709_ _2335_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6118__A2 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6689_ _3241_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7166__I1 mod.Data_Mem.F_M.MRAM\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4129__A1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__C _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8428_ _0524_ net87 mod.Data_Mem.F_M.MRAM\[791\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8359_ _0455_ net226 mod.Data_Mem.F_M.MRAM\[781\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5515__I _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6054__A1 _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A1 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__I mod.Data_Mem.F_M.MRAM\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5425__I _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4540__A1 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5361__S _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7640__I mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4040_ mod.Arithmetic.I_out\[73\] _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout370_I net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5891__I1 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _2524_ _2148_ _2603_ _2605_ _2609_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_92_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7730_ mod.Data_Mem.F_M.MRAM\[795\]\[1\] _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8027__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7661_ _3824_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4873_ _1541_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6612_ _3196_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4359__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7592_ _3604_ _3446_ _3758_ _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8177__CLK net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5020__A2 mod.Data_Mem.F_M.MRAM\[787\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6543_ _2641_ mod.Data_Mem.F_M.MRAM\[769\]\[6\] _2101_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7148__I1 mod.Data_Mem.F_M.MRAM\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ _3003_ _2300_ _3004_ _2512_ _2518_ _3005_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5859__A1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8213_ _0314_ net145 mod.Data_Mem.F_M.MRAM\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5425_ _2079_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6520__A2 mod.Data_Mem.F_M.MRAM\[781\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5356_ _2018_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8144_ mod.Data_Mem.F_M.out_data\[54\] net63 net363 mod.Arithmetic.CN.I_in\[54\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _0894_ _0832_ _0893_ mod.Arithmetic.CN.I_in\[33\] _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8075_ mod.P3.Res\[3\] net32 net245 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5287_ _1931_ _1935_ _1950_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7550__I _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7320__I1 mod.Data_Mem.F_M.MRAM\[770\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5087__A2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7026_ _3248_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5331__I0 mod.Data_Mem.F_M.MRAM\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ _0671_ _0848_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_75_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6166__I _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4169_ _0662_ _0844_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6036__A1 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6036__B2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4598__A1 mod.Arithmetic.ACTI.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7928_ _0154_ net303 mod.Data_Mem.F_M.MRAM\[8\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7859_ _3913_ _3917_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7139__I1 mod.Data_Mem.F_M.MRAM\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4770__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6275__A1 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5078__A2 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5322__I0 mod.Data_Mem.F_M.MRAM\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__I _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A1 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__C _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6502__A2 mod.Data_Mem.F_M.MRAM\[768\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5210_ mod.Data_Mem.F_M.MRAM\[5\]\[4\] mod.Data_Mem.F_M.MRAM\[4\]\[4\] _1874_ _1875_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6190_ _2757_ _2803_ _2804_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4994__I _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5141_ _1761_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5313__I0 mod.Data_Mem.F_M.MRAM\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _1737_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4023_ _0685_ mod.Arithmetic.I_out\[77\] _0695_ _0698_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_96_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4292__A3 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ mod.Data_Mem.F_M.MRAM\[770\]\[5\] mod.Data_Mem.F_M.MRAM\[771\]\[5\] _2490_
+ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7713_ _3850_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout31_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4925_ _1492_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7746__S _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7644_ mod.Data_Mem.F_M.MRAM\[788\]\[6\] _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5529__B1 mod.Data_Mem.F_M.MRAM\[799\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4856_ _1524_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7575_ _3775_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4787_ _0624_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6526_ _2203_ _2327_ _3059_ _2597_ _2598_ _3058_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6457_ mod.Data_Mem.F_M.MRAM\[13\]\[2\] _2375_ _3063_ mod.Data_Mem.F_M.MRAM\[1\]\[2\]
+ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5065__I _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ _1727_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6388_ mod.Data_Mem.F_M.MRAM\[781\]\[7\] _2900_ _2901_ mod.Data_Mem.F_M.MRAM\[780\]\[7\]
+ _2997_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_88_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8127_ mod.Data_Mem.F_M.out_data\[37\] net37 net273 mod.Arithmetic.CN.I_in\[37\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ mod.Data_Mem.F_M.MRAM\[773\]\[6\] mod.Data_Mem.F_M.MRAM\[772\]\[6\] _1908_
+ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8058_ _0267_ net184 mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7009_ _3405_ mod.Data_Mem.F_M.MRAM\[17\]\[7\] _3440_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_169_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6009__A1 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8342__CLK net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6804__I0 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A3 _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6032__I1 mod.Data_Mem.F_M.MRAM\[771\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4043__I0 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7780__I1 mod.Data_Mem.F_M.MRAM\[797\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4080__S _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__A1 mod.Arithmetic.CN.I_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7048__I0 _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5471__A2 mod.Data_Mem.F_M.MRAM\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5859__B _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__B1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6420__A1 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout333_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4710_ _1372_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5690_ _2318_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4641_ _0701_ _0685_ _1061_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7365__I mod.Data_Mem.F_M.MRAM\[772\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5086__S _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5377__I3 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7771__I1 mod.Data_Mem.F_M.MRAM\[797\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7360_ _3653_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4572_ mod.Arithmetic.CN.I_in\[67\] _1128_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6311_ _1577_ _1952_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7291_ _1719_ _3609_ _3611_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8215__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6487__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6242_ _2128_ mod.Data_Mem.F_M.MRAM\[783\]\[3\] mod.Data_Mem.F_M.MRAM\[782\]\[3\]
+ _2064_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6487__B2 _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6173_ _2192_ _2675_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5124_ _1706_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout79_I net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5055_ _1703_ _1709_ _1716_ _1722_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4006_ mod.Arithmetic.I_out\[79\] _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6444__I _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5957_ _1628_ _2141_ _2143_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__S _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _1576_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4973__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ _2158_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7211__I0 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4899__I _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7627_ _3807_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4839_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7275__I mod.Data_Mem.F_M.MRAM\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5922__B1 _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _3308_ _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6112__C _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _3083_ _3102_ _3105_ _3110_ _3113_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_88_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__B _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7489_ _3638_ mod.Data_Mem.F_M.MRAM\[781\]\[1\] _3720_ _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5523__I _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_405 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_416 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_427 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_438 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_449 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5453__A2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3978__I _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6402__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__B _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__B1 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4192__A2 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7505__I1 mod.Data_Mem.F_M.MRAM\[781\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5861__C _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5819__I1 mod.Data_Mem.F_M.MRAM\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout283_I net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__I1 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _3352_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ _2434_ mod.Data_Mem.F_M.MRAM\[773\]\[1\] _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ mod.Data_Mem.F_M.MRAM\[799\]\[3\] _3309_ _3300_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8530_ _0034_ net288 mod.Data_Mem.F_M.out_data\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5742_ _2366_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8461_ _0557_ net157 mod.Data_Mem.F_M.MRAM\[795\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6157__B1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5673_ _2207_ mod.Data_Mem.F_M.MRAM\[797\]\[3\] _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7412_ _3679_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4624_ mod.Arithmetic.CN.I_in\[13\] _1189_ _0971_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8392_ _0488_ net179 mod.Data_Mem.F_M.MRAM\[786\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7343_ _3644_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5380__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4555_ _1226_ _0995_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7274_ _3599_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4486_ _1153_ _1155_ _1156_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_131_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5132__A1 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ _2834_ _2838_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__A2 mod.Data_Mem.F_M.MRAM\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _1568_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5107_ _1706_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _2699_ _2702_ _2703_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_79_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ _1542_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3997__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6989_ _3405_ mod.Data_Mem.F_M.MRAM\[16\]\[7\] _3428_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6902__I _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4410__A3 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7499__I0 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput8 net8 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput10 net10 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5123__A1 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A3 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5202__B _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6084__I _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A1 mod.Data_Mem.F_M.MRAM\[790\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6812__I mod.Data_Mem.F_M.MRAM\[789\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4401__A3 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5428__I _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout129_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5591__C _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4340_ _1009_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_113_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5114__A1 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4271_ _0943_ _0937_ _0944_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5665__A2 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _2345_ _2628_ _2347_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4468__A3 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__A2 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7961_ _0187_ net197 mod.Data_Mem.F_M.MRAM\[779\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6208__B _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6912_ _3249_ mod.Data_Mem.F_M.MRAM\[13\]\[4\] _3381_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7892_ _0118_ net171 mod.Data_Mem.F_M.MRAM\[25\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6217__I1 mod.Data_Mem.F_M.MRAM\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4640__A3 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _3316_ _3337_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6774_ _3295_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3986_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8513_ _0017_ net330 mod.Data_Mem.F_M.out_data\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _2349_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8444_ _0540_ net192 mod.Data_Mem.F_M.MRAM\[793\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5656_ _2284_ _2285_ _2286_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5353__A1 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4607_ _1159_ _1196_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8375_ _0471_ net119 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7553__I _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5587_ _1510_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7326_ _3620_ mod.Data_Mem.F_M.MRAM\[770\]\[7\] _3625_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4538_ _0664_ mod.Arithmetic.CN.I_in\[44\] _0897_ _0983_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_85_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5105__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7257_ mod.Data_Mem.F_M.MRAM\[31\]\[4\] _3312_ _3590_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4469_ _1087_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_77_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6208_ _1737_ _1795_ _2782_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7188_ _3549_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _1804_ _1640_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4417__I mod.Arithmetic.CN.I_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8083__CLK net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4395__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4152__I _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7920__CLK net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5344__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7463__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3991__I _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4698__A3 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6079__I _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5647__A2 mod.Data_Mem.F_M.MRAM\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__A1 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5711__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6743__S _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8576__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5359__S _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout246_I net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4386__A2 mod.Arithmetic.CN.I_in\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7574__S _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5510_ _2136_ mod.Data_Mem.F_M.MRAM\[798\]\[7\] _2151_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6490_ _3082_ _3095_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4138__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5441_ _1553_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4689__A3 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8160_ mod.Data_Mem.F_M.out_data\[70\] net64 net383 mod.Arithmetic.CN.I_in\[70\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5886__A2 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5372_ mod.Data_Mem.F_M.MRAM\[783\]\[7\] _1679_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7111_ _3503_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4323_ _0649_ mod.Arithmetic.CN.I_in\[51\] _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8091_ mod.Data_Mem.F_M.out_data\[1\] net58 net345 mod.Arithmetic.ACTI.x\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout107 net108 net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout118 net119 net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5638__A2 mod.Data_Mem.F_M.MRAM\[797\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ _3467_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout129 net130 net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4254_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5621__I _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4185_ _0754_ _0860_ _0800_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout61_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7944_ _0170_ net190 mod.Data_Mem.F_M.MRAM\[789\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7875_ _0101_ net156 mod.Data_Mem.F_M.MRAM\[24\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6452__I _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ _3271_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5949__I0 mod.Data_Mem.F_M.MRAM\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7943__CLK net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6757_ _3285_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5574__A1 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4377__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3969_ _0639_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5708_ _2077_ _2331_ _2334_ _2302_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6688_ _3240_ mod.Data_Mem.F_M.MRAM\[28\]\[1\] _3237_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7315__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8427_ _0523_ net138 mod.Data_Mem.F_M.MRAM\[791\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5639_ _1706_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8358_ _0454_ net222 mod.Data_Mem.F_M.MRAM\[781\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7309_ _3622_ _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8289_ _0385_ net184 mod.Data_Mem.F_M.MRAM\[772\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8449__CLK net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7626__I0 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5687__B _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__I _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A2 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7193__I _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout196_I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5441__I _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _2454_ _2607_ _2608_ _2529_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_64_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__I0 mod.Data_Mem.F_M.MRAM\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7660_ mod.Data_Mem.F_M.MRAM\[790\]\[6\] _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4872_ mod.Data_Mem.F_M.src\[0\] _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6611_ mod.Data_Mem.F_M.MRAM\[24\]\[1\] _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7591_ _3785_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6542_ _3084_ mod.Data_Mem.F_M.MRAM\[768\]\[6\] _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6473_ _2535_ _3074_ _3078_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8212_ _0313_ net144 mod.Data_Mem.F_M.MRAM\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5424_ mod.Data_Mem.F_M.src\[8\] _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8143_ mod.Data_Mem.F_M.out_data\[53\] net63 net356 mod.Arithmetic.CN.I_in\[53\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5355_ _1998_ _2017_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_99_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4306_ _0644_ mod.Arithmetic.CN.I_in\[35\] _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8074_ mod.P3.Res\[2\] net36 net284 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5286_ _1671_ _1943_ _1949_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7025_ _3455_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4237_ _0670_ _0848_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5331__I1 mod.Data_Mem.F_M.MRAM\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4295__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ _0617_ mod.Arithmetic.CN.I_in\[57\] _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6036__A2 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4099_ _0769_ _0770_ _0754_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6587__A3 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7927_ _0153_ net372 mod.Data_Mem.F_M.MRAM\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7858_ _3931_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6809_ _3323_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5547__A1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8121__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5547__B2 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7789_ _3892_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5727__S _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__I _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6275__A2 _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5322__I1 mod.Data_Mem.F_M.MRAM\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4286__A1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A2 mod.Data_Mem.F_M.MRAM\[786\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7188__I _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6092__I _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6820__I mod.Data_Mem.F_M.MRAM\[789\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__A1 mod.Arithmetic.CN.I_in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout111_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout209_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5710__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5140_ _1674_ _1627_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4496__B _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5071_ mod.Data_Mem.F_M.MRAM\[1\]\[2\] mod.Data_Mem.F_M.MRAM\[0\]\[2\] _1519_ _1738_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5313__I1 mod.Data_Mem.F_M.MRAM\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4022_ _0696_ _0697_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4029__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5077__I0 mod.Data_Mem.F_M.MRAM\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5777__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ _2387_ _2589_ _2592_ _2390_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7712_ mod.Data_Mem.F_M.MRAM\[794\]\[0\] _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4924_ _1587_ _1592_ _1561_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout24_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7643_ _3815_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5529__A1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _1505_ _1523_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5529__B2 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8294__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7574_ _3747_ mod.Data_Mem.F_M.MRAM\[785\]\[1\] _3773_ _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4786_ mod.Arithmetic.CN.I_in\[15\] _1455_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4201__A1 mod.Arithmetic.CN.I_in\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6525_ _2548_ _2589_ _3124_ _3125_ _3128_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ _2498_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5407_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6387_ _2902_ _2996_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8126_ mod.Data_Mem.F_M.out_data\[36\] net30 net273 mod.Arithmetic.CN.I_in\[36\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5338_ mod.Data_Mem.F_M.MRAM\[771\]\[6\] mod.Data_Mem.F_M.MRAM\[770\]\[6\] _1906_
+ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8057_ _0266_ net147 mod.Data_Mem.F_M.MRAM\[20\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6501__I0 mod.Data_Mem.F_M.MRAM\[780\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5269_ _1933_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7008_ _3443_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6009__A2 mod.Data_Mem.F_M.MRAM\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6804__I1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6841__S _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4440__A1 mod.Arithmetic.CN.I_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6193__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4043__I1 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5240__I0 mod.Data_Mem.F_M.MRAM\[773\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5940__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5256__I _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__A2 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__S0 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8174__RN net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6248__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4259__A1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8167__CLK net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout290 net295 net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_93_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7048__I1 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__B2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout159_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4431__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5367__S _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7646__I mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4640_ _0614_ mod.Arithmetic.CN.I_in\[22\] _0684_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout326_I net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5931__A1 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ mod.Arithmetic.CN.I_in\[66\] _1129_ _0648_ _0781_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7582__S _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6310_ _2893_ _2920_ _2921_ _2881_ _2072_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7290_ _3610_ _3609_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8165__RN net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6241_ _1637_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6487__A2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7381__I mod.Data_Mem.F_M.MRAM\[773\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6172_ _2743_ _2752_ _2787_ _2367_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_44_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5123_ _1786_ mod.Data_Mem.F_M.MRAM\[789\]\[2\] _1789_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6926__S _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _1602_ _1721_ _1617_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4005_ _0680_ mod.Arithmetic.I_out\[79\] _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4670__A1 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5956_ _2548_ _2572_ _2575_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4422__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4907_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5887_ _2117_ _2494_ _2508_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5277__S _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7211__I1 mod.Data_Mem.F_M.MRAM\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7626_ _3806_ mod.Data_Mem.F_M.MRAM\[787\]\[5\] _3801_ _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4838_ _1500_ _1506_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6175__A1 _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7557_ _1797_ _3762_ _3764_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5922__A1 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _0624_ _1134_ mod.Arithmetic.CN.I_in\[61\] _1366_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5922__B2 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6508_ _1491_ _3112_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5009__C _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7488_ _3721_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6439_ _2090_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8109_ mod.Data_Mem.F_M.out_data\[19\] net46 net329 mod.Arithmetic.CN.I_in\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_406 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_417 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_428 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_439 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6402__A2 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4413__A1 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__I0 mod.Data_Mem.F_M.MRAM\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__I0 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5913__B2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5915__S _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6469__A2 mod.Data_Mem.F_M.MRAM\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8147__RN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6713__I0 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6746__S _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout276_I net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _2224_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6790_ _3308_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _1547_ _1532_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5097__S _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6280__I _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8460_ _0556_ net173 mod.Data_Mem.F_M.MRAM\[795\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5672_ _2131_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6157__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6157__B2 _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7411_ mod.Data_Mem.F_M.MRAM\[775\]\[6\] _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4623_ _1292_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8391_ _0487_ net77 mod.Data_Mem.F_M.MRAM\[785\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6952__I0 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5825__S _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7342_ _3615_ mod.Data_Mem.F_M.MRAM\[771\]\[4\] _3643_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4554_ mod.Arithmetic.CN.I_in\[52\] _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5380__A2 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4949__B _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8332__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8138__RN net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7273_ mod.Data_Mem.F_M.MRAM\[5\]\[4\] _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4485_ _1087_ _1141_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout91_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6224_ mod.Data_Mem.F_M.MRAM\[13\]\[3\] _2193_ _2836_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6155_ _2701_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5106_ _1662_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _1830_ _1616_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ mod.Data_Mem.F_M.MRAM\[773\]\[1\] mod.Data_Mem.F_M.MRAM\[772\]\[1\] _1704_
+ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4643__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7487__S _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6988_ _3431_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5939_ _2136_ mod.Data_Mem.F_M.MRAM\[3\]\[4\] _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_107_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7609_ _3784_ mod.Data_Mem.F_M.MRAM\[786\]\[7\] _3786_ _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8589_ _0605_ net167 mod.Data_Mem.F_M.MRAM\[9\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8129__RN net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7499__I1 mod.Data_Mem.F_M.MRAM\[781\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput9 net9 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5534__I _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5123__A2 mod.Data_Mem.F_M.MRAM\[789\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4882__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7120__I0 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7820__A1 _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4634__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5202__C _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4937__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7196__I _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A1 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _0867_ _0936_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6311__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5114__A2 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout393_I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7960_ _0186_ net161 mod.Data_Mem.F_M.MRAM\[779\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6911_ _3375_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7891_ _0117_ net173 mod.Data_Mem.F_M.MRAM\[25\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6217__I2 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _3343_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6378__A1 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4951__C _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6773_ mod.Data_Mem.F_M.dest\[1\] mod.Data_Mem.F_M.dest\[0\] _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3985_ _0661_ mod.Arithmetic.CN.I_in\[56\] _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5619__I _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__I _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5724_ _2166_ _1500_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8512_ _0016_ net340 mod.Data_Mem.F_M.out_data\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8443_ _0539_ net166 mod.Data_Mem.F_M.MRAM\[793\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5655_ _2264_ _2124_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4606_ _1154_ _1275_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8374_ _0470_ net119 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6550__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5586_ _1580_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4156__A3 mod.Arithmetic.CN.I_in\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7325_ _3632_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4537_ _0659_ _1208_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7256_ _3584_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6302__A1 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5105__A2 mod.Data_Mem.F_M.MRAM\[771\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4468_ _1103_ _1108_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6207_ _2774_ _1799_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7187_ _3294_ _3464_ _3335_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_58_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4399_ _1068_ _1069_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6138_ _2325_ mod.Data_Mem.F_M.MRAM\[6\]\[1\] mod.Data_Mem.F_M.MRAM\[7\]\[1\] _2753_
+ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ mod.Data_Mem.F_M.MRAM\[781\]\[0\] _2685_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8228__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7169__I0 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6916__I0 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6541__A1 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5344__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6844__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4855__A1 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5439__I _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5032__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout141_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout239_I net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6907__I0 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__S _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5335__A2 _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6532__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5371_ _2019_ _2025_ _2026_ _2032_ _1900_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7590__S _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7110_ _3450_ mod.Data_Mem.F_M.MRAM\[3\]\[1\] _3501_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4322_ _0658_ mod.Arithmetic.CN.I_in\[50\] _0842_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8090_ mod.Data_Mem.F_M.out_data\[0\] net54 net344 mod.Arithmetic.ACTI.x\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout108 net112 net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7041_ _3445_ mod.Data_Mem.F_M.MRAM\[1\]\[0\] _3466_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout119 net120 net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4253_ mod.Arithmetic.CN.I_in\[50\] _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5902__I _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4184_ _0769_ _0770_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout54_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7943_ _0169_ net154 mod.Data_Mem.F_M.MRAM\[789\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5271__A1 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7874_ _0100_ net172 mod.Data_Mem.F_M.MRAM\[24\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6825_ _3331_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5949__I1 mod.Data_Mem.F_M.MRAM\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5023__A1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7765__S _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6756_ mod.Data_Mem.F_M.MRAM\[8\]\[1\] _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5574__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3968_ _0644_ mod.Arithmetic.CN.I_in\[16\] _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5707_ _2277_ _2148_ _2332_ _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6687_ _3239_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8426_ _0522_ net188 mod.Data_Mem.F_M.MRAM\[791\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6523__A1 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5638_ _2269_ mod.Data_Mem.F_M.MRAM\[797\]\[1\] _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5731__C1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8357_ _0453_ net230 mod.Data_Mem.F_M.MRAM\[781\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5569_ _2054_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7308_ _3332_ _3604_ _3446_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8288_ _0384_ net150 mod.Data_Mem.F_M.MRAM\[772\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7239_ _3580_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7005__S _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4837__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4301__A3 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7626__I1 mod.Data_Mem.F_M.MRAM\[787\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A3 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A2 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5262__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6514__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5317__A2 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6818__I mod.Data_Mem.F_M.MRAM\[789\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout189_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4940_ _1541_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout356_I net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4851__I1 mod.Data_Mem.F_M.MRAM\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ _1529_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ _3195_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7590_ _3784_ mod.Data_Mem.F_M.MRAM\[785\]\[7\] _3779_ _3785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6541_ _2089_ _2613_ _3143_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6472_ _3020_ _2517_ _2513_ _3004_ _3077_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6505__A1 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__B2 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8211_ _0312_ net161 mod.Data_Mem.F_M.MRAM\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5423_ _2078_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6929__S _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8073__CLK net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5354_ _1999_ _2005_ _2016_ _1931_ _1630_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8142_ mod.Data_Mem.F_M.out_data\[52\] net63 net354 mod.Arithmetic.CN.I_in\[52\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6269__B1 _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4305_ _0896_ _0900_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8073_ mod.P3.Res\[1\] net32 net246 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5285_ _1808_ _1946_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7024_ _3454_ mod.Data_Mem.F_M.MRAM\[18\]\[3\] _3448_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4236_ _0845_ _0909_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4295__A2 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5492__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4167_ _0660_ _0842_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_110_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7910__CLK net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4098_ _0760_ _0772_ _0773_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7926_ _0152_ net157 mod.Data_Mem.F_M.MRAM\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7857_ mod.Data_Mem.F_M.MRAM\[9\]\[7\] _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5079__I _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6808_ mod.Data_Mem.F_M.MRAM\[799\]\[7\] _3322_ _3313_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5547__A2 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7788_ _3306_ mod.Data_Mem.F_M.MRAM\[798\]\[2\] _3889_ _3892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4755__B1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6739_ _3240_ mod.Data_Mem.F_M.MRAM\[0\]\[1\] _3274_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5807__I _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7544__I0 _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8409_ _0505_ net160 mod.Data_Mem.F_M.MRAM\[788\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4507__B1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6839__S _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4286__A2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5483__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4158__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5235__A1 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8505__D _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A3 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6735__A1 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout90 net93 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4210__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8096__CLK net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout104_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5710__A2 mod.Data_Mem.F_M.MRAM\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__C _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7933__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ _1732_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4021_ _0696_ _0697_ _0686_ _0687_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_81_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7379__I mod.Data_Mem.F_M.MRAM\[773\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__I1 mod.Data_Mem.F_M.MRAM\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__B1 _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6423__C2 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5972_ _2590_ mod.Data_Mem.F_M.MRAM\[772\]\[5\] _2591_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5777__A2 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7711_ _3849_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ _1589_ _1590_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6026__I0 mod.Data_Mem.F_M.MRAM\[784\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7642_ mod.Data_Mem.F_M.MRAM\[788\]\[5\] _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4854_ _1522_ _1492_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5529__A2 mod.Data_Mem.F_M.MRAM\[798\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7774__I0 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout17_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4785_ _1289_ _0737_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6232__B _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7573_ _3774_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4201__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4531__I _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ _2488_ _2594_ _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _2861_ _3053_ _3061_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5406_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6386_ _2268_ mod.Data_Mem.F_M.MRAM\[783\]\[7\] mod.Data_Mem.F_M.MRAM\[782\]\[7\]
+ _2904_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5337_ mod.Data_Mem.F_M.MRAM\[769\]\[6\] mod.Data_Mem.F_M.MRAM\[768\]\[6\] _1904_
+ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8125_ mod.Data_Mem.F_M.out_data\[35\] net47 net278 mod.Arithmetic.CN.I_in\[35\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5268_ _1901_ _1932_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_60_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8056_ _0265_ net147 mod.Data_Mem.F_M.MRAM\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6501__I1 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7007_ _3403_ mod.Data_Mem.F_M.MRAM\[17\]\[6\] _3440_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4219_ mod.Arithmetic.CN.I_in\[34\] _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _1489_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5768__A2 mod.Data_Mem.F_M.MRAM\[788\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7909_ _0135_ net236 mod.Data_Mem.F_M.MRAM\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6017__I0 mod.Data_Mem.F_M.MRAM\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4440__A2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7765__I0 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5537__I _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__A2 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8194__574 net574 vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5940__A2 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5379__S1 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5473__S _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7956__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5272__I _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4259__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout280 net281 net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout291 net294 net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5759__A2 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6036__C _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__I _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5875__C _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout221_I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4195__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout319_I net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4570_ _0667_ mod.Arithmetic.CN.I_in\[69\] _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5931__A2 mod.Data_Mem.F_M.MRAM\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6240_ mod.Data_Mem.F_M.MRAM\[781\]\[3\] _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6171_ _2219_ _2770_ _2778_ _2786_ _2737_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5122_ _1787_ _1788_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5115__C _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5447__A1 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5053_ _1717_ mod.Data_Mem.F_M.MRAM\[769\]\[1\] _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4004_ mod.Arithmetic.CN.I_in\[15\] _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5955_ _2390_ _2573_ _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _1574_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5886_ _2372_ _2497_ _2507_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_33_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7625_ _3315_ _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4837_ _1502_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7556_ _3612_ _3762_ _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ mod.Arithmetic.ACTI.x\[7\] _1436_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6507_ _3049_ _3111_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4699_ _0658_ mod.Arithmetic.CN.I_in\[69\] _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7487_ _3718_ mod.Data_Mem.F_M.MRAM\[781\]\[0\] _3720_ _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6438_ _3026_ _2442_ _3045_ _3005_ _1623_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6369_ _2027_ _2028_ _1746_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8108_ mod.Data_Mem.F_M.out_data\[18\] net54 net349 mod.Arithmetic.CN.I_in\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_407 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8039_ _0248_ net191 mod.Data_Mem.F_M.MRAM\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtiny_user_project_418 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_429 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5820__I _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4661__A2 mod.Arithmetic.CN.I_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8092__RN net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4413__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5610__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5610__B2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5461__I1 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A2 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6961__I1 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6713__I1 mod.Data_Mem.F_M.MRAM\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8134__CLK net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5677__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A1 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5730__I _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6492__I3 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout171_I net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout269_I net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5601__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4404__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5740_ _2346_ _2356_ _2364_ _1499_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5671_ _2070_ _2300_ _2162_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6157__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4081__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7410_ _3678_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4168__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4622_ _0737_ _1191_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8390_ _0486_ net74 mod.Data_Mem.F_M.MRAM\[785\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__I1 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7341_ _3635_ _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4553_ _1118_ _1119_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5905__I _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7272_ _3598_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4484_ _1087_ _1141_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5668__A1 _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6223_ _1622_ _2695_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _2761_ _2769_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout84_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__I _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5105_ _1767_ mod.Data_Mem.F_M.MRAM\[771\]\[2\] _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6085_ _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5036_ _1609_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4643__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6987_ _3403_ mod.Data_Mem.F_M.MRAM\[16\]\[6\] _3428_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8074__RN net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5288__S _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8007__CLK net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _2100_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ mod.Data_Mem.F_M.MRAM\[784\]\[3\] mod.Data_Mem.F_M.MRAM\[785\]\[3\] _2490_
+ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7608_ _3795_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8588_ _0604_ net197 mod.Data_Mem.F_M.MRAM\[9\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7539_ _3725_ _1902_ _3752_ _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5659__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6847__S _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8527__562 net562 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4882__A2 _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5550__I _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4634__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A1 mod.Arithmetic.CN.I_in\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5595__B1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5725__I _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4570__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6311__A2 _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4322__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout386_I net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6075__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5822__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6910_ _3380_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7890_ _0116_ net170 mod.Data_Mem.F_M.MRAM\[25\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _3249_ mod.Data_Mem.F_M.MRAM\[769\]\[4\] _3340_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6217__I3 mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6291__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _3229_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3984_ _0616_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6224__C _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8511_ net570 net358 mod.Data_Mem.F_M.out_data\[71\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5723_ _2347_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8442_ _0538_ net156 mod.Data_Mem.F_M.MRAM\[793\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5654_ _2271_ mod.Data_Mem.F_M.MRAM\[796\]\[2\] _2262_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4605_ _1158_ _1259_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4936__I0 mod.Data_Mem.F_M.MRAM\[789\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8373_ _0469_ net127 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6550__A2 mod.Data_Mem.F_M.MRAM\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ _1599_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7324_ _3618_ mod.Data_Mem.F_M.MRAM\[770\]\[6\] _3625_ _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4536_ mod.Arithmetic.CN.I_in\[45\] _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _3589_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4467_ _1121_ _1122_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_85_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ _1608_ _1790_ _2733_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4313__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7186_ _3548_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4398_ mod.Arithmetic.CN.I_in\[26\] _1064_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _2225_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A1 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6068_ _2684_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5813__A1 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__B2 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5019_ _1515_ _1686_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__B1 mod.Data_Mem.F_M.MRAM\[798\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7318__A1 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7169__I1 mod.Data_Mem.F_M.MRAM\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6526__C1 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6916__I1 mod.Data_Mem.F_M.MRAM\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4552__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4304__B2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4855__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5804__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7201__S _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7557__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5032__A2 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5583__A3 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__A1 mod.Arithmetic.CN.I_in\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout134_I net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__C1 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6907__I1 mod.Data_Mem.F_M.MRAM\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6532__A2 mod.Data_Mem.F_M.MRAM\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout301_I net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _1671_ _2031_ _1624_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4321_ _0658_ _0928_ mod.Arithmetic.CN.I_in\[51\] _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_114_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6296__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7040_ _3465_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout109 net111 net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4252_ _0911_ _0921_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_99_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4183_ _0858_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ _0168_ net138 mod.Data_Mem.F_M.MRAM\[789\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7873_ _0099_ net316 mod.Data_Mem.F_M.MRAM\[24\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout47_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ mod.Data_Mem.F_M.MRAM\[789\]\[7\] _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5023__A2 mod.Data_Mem.F_M.MRAM\[789\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6220__A1 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ _3284_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3967_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ _2315_ mod.Data_Mem.F_M.MRAM\[796\]\[6\] _2280_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ net4 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8425_ _0521_ net150 mod.Data_Mem.F_M.MRAM\[791\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5637_ _2268_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6523__A2 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5731__B1 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8356_ _0452_ net221 mod.Data_Mem.F_M.MRAM\[781\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5568_ mod.Data_Mem.F_M.MRAM\[29\]\[3\] _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5731__C2 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7307_ _3621_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4519_ _0730_ _0713_ _0971_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8287_ _0383_ net121 mod.Data_Mem.F_M.MRAM\[771\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5499_ _2142_ mod.Data_Mem.F_M.MRAM\[31\]\[5\] _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238_ _3533_ mod.Data_Mem.F_M.MRAM\[30\]\[4\] _3579_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4837__A2 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7169_ _3539_ mod.Data_Mem.F_M.MRAM\[12\]\[7\] _3534_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8524__565 net565 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6834__I0 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7021__S _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8495__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5476__S _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6514__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6278__A1 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5325__I0 mod.Data_Mem.F_M.MRAM\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout251_I net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout349_I net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4870_ _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6202__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7250__I0 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7862__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6540_ _2611_ mod.Data_Mem.F_M.MRAM\[780\]\[6\] _3142_ _2168_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4764__B2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6471_ _2414_ _3075_ _3076_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_9_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6505__A2 _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ _0311_ net243 mod.Data_Mem.F_M.MRAM\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4516__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5422_ _1805_ _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8141_ mod.Data_Mem.F_M.out_data\[51\] net55 net354 mod.Arithmetic.CN.I_in\[51\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5353_ mod.Data_Mem.F_M.MRAM\[799\]\[6\] _1914_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6269__A1 _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6269__B2 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4304_ _0902_ _0903_ _0934_ _0977_ _0908_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__5316__I0 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8072_ mod.P3.Res\[0\] net61 net384 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5284_ _1569_ _1947_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4819__A2 _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7023_ _3245_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4235_ _0655_ _0665_ mod.Arithmetic.CN.I_in\[64\] _0849_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_101_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5492__A2 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4166_ _0617_ mod.Arithmetic.CN.I_in\[49\] _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4097_ mod.Arithmetic.ACTI.x\[2\] _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7925_ _0151_ net125 mod.Data_Mem.F_M.MRAM\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6992__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7856_ _3930_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6807_ _3321_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7787_ _3891_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4999_ mod.Data_Mem.F_M.MRAM\[22\]\[1\] _1643_ _1666_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4755__A1 mod.Arithmetic.CN.I_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6738_ _3275_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4755__B2 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ mod.Data_Mem.F_M.MRAM\[27\]\[6\] _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5095__I _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7544__I1 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4507__A1 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8408_ _0504_ net140 mod.Data_Mem.F_M.MRAM\[788\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8339_ _0435_ net308 mod.Data_Mem.F_M.MRAM\[778\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5823__I _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5483__A2 mod.Data_Mem.F_M.MRAM\[798\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A1 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7480__I0 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6283__I1 _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8521__D _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4746__A1 mod.Arithmetic.CN.I_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout80 net84 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout91 net93 net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6499__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5171__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8510__CLK net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout299_I net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4020_ mod.Arithmetic.CN.I_in\[20\] _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5474__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6423__A1 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__B2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5971_ _2351_ mod.Data_Mem.F_M.MRAM\[773\]\[5\] _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_92_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7710_ mod.Data_Mem.F_M.MRAM\[793\]\[7\] _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4922_ _1564_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7223__I0 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7641_ _3814_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4037__I0 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4853_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7774__I1 mod.Data_Mem.F_M.MRAM\[797\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5908__I _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7572_ _3771_ mod.Data_Mem.F_M.MRAM\[785\]\[0\] _3773_ _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4784_ _0744_ _1295_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _2632_ _1955_ _2399_ _3126_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5844__S _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6454_ _3054_ _3055_ _3060_ _3013_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8190__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6385_ mod.Data_Mem.F_M.MRAM\[13\]\[7\] _1538_ _2194_ mod.Data_Mem.F_M.MRAM\[12\]\[7\]
+ _2994_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_88_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8124_ mod.Data_Mem.F_M.out_data\[34\] net59 net355 mod.Arithmetic.CN.I_in\[34\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5336_ mod.Data_Mem.F_M.MRAM\[783\]\[6\] _1702_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8055_ _0264_ net163 mod.Data_Mem.F_M.MRAM\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6111__B1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5267_ _1903_ _1913_ _1930_ _1931_ _1630_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6501__I2 mod.Data_Mem.F_M.MRAM\[781\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7006_ _3442_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5465__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4218_ _0644_ mod.Arithmetic.CN.I_in\[34\] _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5198_ mod.Data_Mem.F_M.MRAM\[783\]\[3\] _1863_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4149_ _0621_ _0656_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7908_ _0134_ net242 mod.Data_Mem.F_M.MRAM\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__I1 mod.Data_Mem.F_M.MRAM\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7839_ _3169_ _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7765__I1 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8533__CLK net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5153__A1 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4259__A3 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout270 net271 net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout281 net282 net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout292 net294 net292 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6405__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7205__I0 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5728__I _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__I _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4719__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout214_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6170_ _1807_ _2785_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5121_ mod.Data_Mem.F_M.MRAM\[788\]\[2\] _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5447__A2 mod.Data_Mem.F_M.MRAM\[799\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5052_ _1718_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4003_ mod.Arithmetic.CN.I_in\[23\] _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4958__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5954_ _2391_ mod.Data_Mem.F_M.MRAM\[20\]\[5\] _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4905_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8556__CLK net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ _2499_ _2502_ _2505_ _2506_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7624_ _1922_ _3804_ _3805_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4836_ _1503_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7555_ _1683_ _3762_ _3763_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5383__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ mod.Arithmetic.CN.I_in\[68\] _1377_ _1422_ mod.Arithmetic.ACTI.x\[5\] _1437_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6506_ _3047_ _2317_ _2488_ _2532_ _2530_ _2559_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7486_ _3719_ _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4698_ _0636_ _1367_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5135__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6437_ mod.Data_Mem.F_M.MRAM\[0\]\[1\] mod.Data_Mem.F_M.MRAM\[1\]\[1\] _2252_ _3045_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6368_ _2867_ _2977_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8107_ mod.Data_Mem.F_M.out_data\[17\] net54 net341 mod.Arithmetic.CN.I_in\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_103_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5319_ _1491_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6299_ _2696_ _2911_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8038_ _0247_ net74 mod.Data_Mem.F_M.MRAM\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtiny_user_project_408 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_419 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A3 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output10_I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5677__A2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6047__C _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4652__A3 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8579__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout164_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _2295_ _2299_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4621_ _0834_ _1290_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4168__A2 mod.Arithmetic.CN.I_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7340_ _3642_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4552_ _0929_ _1113_ _1115_ _1116_ _1112_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5117__A1 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6289__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7271_ mod.Data_Mem.F_M.MRAM\[5\]\[3\] _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4483_ _1047_ _1084_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5668__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _1569_ _2835_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6153_ _2674_ _2764_ _2768_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7114__S _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5104_ _1769_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout77_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6084_ _2700_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6238__B _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7290__A1 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _1565_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6986_ _3430_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5937_ _2434_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7784__S _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _1712_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_167_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7607_ _3782_ mod.Data_Mem.F_M.MRAM\[786\]\[6\] _3786_ _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4819_ _1268_ _1485_ _1486_ _1487_ _1488_ mod.P3.Res\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__4159__A2 mod.Arithmetic.CN.I_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8587_ _0603_ net371 mod.Data_Mem.F_M.MRAM\[9\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5799_ _2415_ _2121_ _2417_ _2396_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_7538_ _3744_ _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_108_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5317__B _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7469_ _3709_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5659__A2 mod.Data_Mem.F_M.MRAM\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7024__S _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5595__A1 mod.Data_Mem.F_M.MRAM\[797\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4398__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5595__B2 mod.Data_Mem.F_M.MRAM\[796\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8101__CLK net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5347__A1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4570__A2 mod.Arithmetic.CN.I_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout281_I net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout379_I net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5822__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6840_ _3342_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6771_ _3292_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3983_ _0659_ mod.Arithmetic.CN.I_in\[48\] _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8510_ net571 net383 mod.Data_Mem.F_M.out_data\[70\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5722_ _2114_ _1534_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8441_ _0537_ net198 mod.Data_Mem.F_M.MRAM\[793\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5653_ _2269_ mod.Data_Mem.F_M.MRAM\[797\]\[2\] _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6521__B _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6535__B1 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4820__I mod.Data_Mem.F_M.src\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _1158_ _1259_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8372_ _0468_ net229 mod.Data_Mem.F_M.MRAM\[783\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5584_ _1554_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4936__I1 mod.Data_Mem.F_M.MRAM\[788\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7323_ _3631_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4535_ _1206_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5852__S _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7254_ mod.Data_Mem.F_M.MRAM\[31\]\[3\] _3555_ _3585_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4466_ _1133_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6205_ _1920_ _1785_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5510__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4313__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ mod.Data_Mem.F_M.MRAM\[22\]\[7\] _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4397_ _0639_ mod.Arithmetic.CN.I_in\[28\] _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _2696_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__A2 _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ _2678_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5018_ mod.Data_Mem.F_M.MRAM\[786\]\[1\] _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5577__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _3419_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7318__A2 _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6526__B1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6526__C2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5501__A1 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__A2 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4068__A1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5804__A2 mod.Data_Mem.F_M.MRAM\[771\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7557__A2 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4240__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6517__B1 _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__C2 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout127_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4543__A2 mod.Arithmetic.CN.I_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5740__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4320_ _0922_ _0663_ _0844_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4251_ _0923_ _0924_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5343__I1 mod.Data_Mem.F_M.MRAM\[788\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4182_ _0803_ mod.P2.Rout_reg\[1\] _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input1_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6453__C1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7941_ _0167_ net98 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8147__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6516__B _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7872_ _0098_ net320 mod.Data_Mem.F_M.MRAM\[24\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _3330_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5559__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6220__A2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6754_ mod.Data_Mem.F_M.MRAM\[8\]\[0\] _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4231__A1 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3966_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5705_ _2128_ mod.Data_Mem.F_M.MRAM\[797\]\[6\] _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6685_ _3238_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5636_ _2053_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8424_ _0520_ net147 mod.Data_Mem.F_M.MRAM\[791\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5031__I0 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8355_ _0451_ net254 mod.Data_Mem.F_M.MRAM\[781\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5731__A1 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5567_ _1600_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7306_ _3620_ mod.Data_Mem.F_M.MRAM\[768\]\[7\] _3608_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4518_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8286_ _0382_ net121 mod.Data_Mem.F_M.MRAM\[771\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5498_ _2053_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7237_ _3573_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6477__I _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4449_ _1007_ _1015_ _1016_ _1105_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_120_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7168_ _3258_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6119_ _2689_ _1498_ _2731_ _2735_ _1865_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7099_ _3496_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5098__I0 mod.Data_Mem.F_M.MRAM\[773\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6834__I1 mod.Data_Mem.F_M.MRAM\[769\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5798__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6426__B _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5757__S _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A2 _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4222__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5556__I _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5722__A1 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5325__I1 mod.Data_Mem.F_M.MRAM\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__S0 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5789__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6450__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7011__I _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6202__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7250__I1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout244_I net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5261__I0 mod.Data_Mem.F_M.MRAM\[785\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A1 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5466__I _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6071__B _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6470_ _2261_ mod.Data_Mem.F_M.MRAM\[12\]\[3\] _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5421_ _2061_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4516__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8195__RN net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5713__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8140_ mod.Data_Mem.F_M.out_data\[50\] net55 net354 mod.Arithmetic.CN.I_in\[50\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5352_ _2007_ _2014_ _1780_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6269__A2 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4303_ _0927_ _0933_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8071_ mod.DMen_reg net25 net237 mod.DMen_reg2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5283_ mod.Data_Mem.F_M.MRAM\[785\]\[5\] mod.Data_Mem.F_M.MRAM\[784\]\[5\] _1874_
+ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7022_ _3453_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4819__A3 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4234_ _0666_ _0849_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _0663_ _0673_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7122__S _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4096_ _0755_ _0714_ _0768_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6246__B _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8164__D mod.Data_Mem.F_M.out_data\[74\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6961__S _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7924_ _0150_ net123 mod.Data_Mem.F_M.MRAM\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4452__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7855_ mod.Data_Mem.F_M.MRAM\[9\]\[6\] _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6806_ net10 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4998_ _1529_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7786_ _3303_ mod.Data_Mem.F_M.MRAM\[798\]\[1\] _3889_ _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6737_ _3228_ mod.Data_Mem.F_M.MRAM\[0\]\[0\] _3274_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3949_ _0626_ mod.DM_en vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4755__A2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _3224_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8407_ _0503_ net97 mod.Data_Mem.F_M.MRAM\[787\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5619_ _1956_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6752__I0 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4507__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__A1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6599_ mod.Data_Mem.F_M.MRAM\[11\]\[3\] _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8338_ _0434_ net375 mod.Data_Mem.F_M.MRAM\[778\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8269_ _0365_ net122 mod.Data_Mem.F_M.MRAM\[768\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8462__CLK net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7480__I1 mod.Data_Mem.F_M.MRAM\[780\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8110__RN net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7766__I _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6196__A1 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5943__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4746__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout70 net76 net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout81 net82 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout92 net93 net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8177__RN net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__I0 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5171__A2 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout194_I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4682__A1 mod.Arithmetic.CN.I_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8101__RN net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6423__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5970_ _1840_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ mod.Data_Mem.F_M.MRAM\[769\]\[0\] mod.Data_Mem.F_M.MRAM\[768\]\[0\] _1585_
+ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4985__A2 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7223__I1 mod.Data_Mem.F_M.MRAM\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7640_ mod.Data_Mem.F_M.MRAM\[788\]\[4\] _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4852_ mod.Data_Mem.F_M.src\[0\] _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6187__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7571_ _3772_ _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4783_ _0743_ _1190_ _1188_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_165_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6522_ _2315_ mod.Data_Mem.F_M.MRAM\[768\]\[5\] _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6453_ _2492_ _2467_ _3057_ _3058_ _3059_ _2466_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7117__S _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5404_ _1594_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _1568_ _2993_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8123_ mod.Data_Mem.F_M.out_data\[33\] net58 net346 mod.Arithmetic.CN.I_in\[33\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5335_ _1984_ _1990_ _1991_ _1997_ _1900_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6956__S _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8054_ _0263_ net125 mod.Data_Mem.F_M.MRAM\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5266_ _1655_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7005_ _3416_ mod.Data_Mem.F_M.MRAM\[17\]\[5\] _3440_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6501__I3 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4217_ _0833_ _0838_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5799__C _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5197_ _1655_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4673__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4148_ mod.Arithmetic.CN.I_in\[32\] _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7611__A1 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4079_ _0716_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__I0 mod.Data_Mem.F_M.MRAM\[798\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _0133_ net235 mod.Data_Mem.F_M.MRAM\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6178__A1 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7838_ _3920_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7769_ _3306_ mod.Data_Mem.F_M.MRAM\[797\]\[2\] _3878_ _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8159__RN net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5689__B1 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5153__A2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout260 net286 net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout271 net272 net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4664__A1 mod.Arithmetic.CN.I_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout282 net283 net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout293 net294 net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6405__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8208__CLK net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4416__A1 _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5613__B1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7496__I _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7205__I1 mod.Data_Mem.F_M.MRAM\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4913__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5216__I0 mod.Data_Mem.F_M.MRAM\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8358__CLK net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6964__I0 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5744__I _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout207_I net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _1609_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7141__I0 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5051_ mod.Data_Mem.F_M.MRAM\[768\]\[1\] _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4002_ mod.Arithmetic.ACTI.x\[7\] _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4095__I _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4407__A1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__B1 mod.Data_Mem.F_M.MRAM\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5953_ _2526_ mod.Data_Mem.F_M.MRAM\[21\]\[5\] _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6524__B _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5919__I _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4823__I mod.Data_Mem.F_M.src\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _1527_ _1545_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5884_ _2115_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout22_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7623_ _3312_ _3804_ _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5907__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4835_ mod.Data_Mem.F_M.src\[1\] _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7554_ _3610_ _3762_ _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5383__A2 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _1422_ mod.Arithmetic.ACTI.x\[7\] _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6505_ _2603_ _2537_ _3106_ _2204_ _3109_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7485_ _3634_ _3371_ _3387_ _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4697_ _1134_ _1251_ _1366_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6436_ _2308_ _2449_ _3043_ _3003_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5135__A2 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6367_ _2973_ _2974_ _2975_ _2976_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5318_ _1965_ _1974_ _1975_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8106_ mod.Data_Mem.F_M.out_data\[16\] net42 net275 mod.Arithmetic.CN.I_in\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_88_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7132__I0 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6298_ _2228_ _2232_ _2907_ _2910_ _2079_ _2744_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8037_ _0246_ net73 mod.Data_Mem.F_M.MRAM\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5249_ _1678_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_409 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4646__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7310__S _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4949__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8500__CLK net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7199__I0 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5564__I _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6323__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6323__B2 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6395__I _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4908__I _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5429__A3 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4844__S _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6344__B _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5062__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout157_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4620_ _0743_ mod.Arithmetic.CN.I_in\[13\] _1190_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout324_I net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6562__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7898__CLK net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4551_ _1121_ _1221_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7106__A3 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7270_ _3597_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6314__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4482_ _0988_ _1083_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _2210_ mod.Data_Mem.F_M.MRAM\[14\]\[3\] mod.Data_Mem.F_M.MRAM\[15\]\[3\] _2278_
+ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _1643_ _2765_ _2766_ _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7114__I0 _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5103_ mod.Data_Mem.F_M.MRAM\[770\]\[2\] _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ _1552_ _1546_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4628__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _1678_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7290__A2 _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5053__A1 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6985_ _3416_ mod.Data_Mem.F_M.MRAM\[16\]\[5\] _3428_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6250__B1 _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _2370_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ mod.Data_Mem.F_M.MRAM\[788\]\[3\] mod.Data_Mem.F_M.MRAM\[789\]\[3\] _2427_
+ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7606_ _3794_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4818_ _0679_ _0680_ mod.Arithmetic.I_out\[79\] _0681_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__6553__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8586_ _0602_ net378 mod.Data_Mem.F_M.MRAM\[9\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5798_ _2418_ _1689_ _2419_ _2421_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7537_ _3751_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4749_ _0623_ mod.Arithmetic.CN.I_in\[70\] _1379_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6305__A1 _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7468_ _3638_ mod.Data_Mem.F_M.MRAM\[780\]\[1\] _3707_ _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6419_ _2618_ _3027_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7399_ mod.Data_Mem.F_M.MRAM\[775\]\[0\] _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8053__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4619__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6943__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6164__B _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5595__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5347__A2 mod.Data_Mem.F_M.MRAM\[786\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7215__S _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4322__A3 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7014__I _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout274_I net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6770_ net3 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3982_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5721_ _2345_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8440_ _0536_ net320 mod.Data_Mem.F_M.MRAM\[793\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6535__A1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _2089_ _1806_ _2276_ _2283_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6535__B2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _0625_ _0738_ _1190_ _1079_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_129_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8371_ _0467_ net255 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5583_ _2219_ _2154_ _2091_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_129_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8076__CLK net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7322_ _3569_ mod.Data_Mem.F_M.MRAM\[770\]\[5\] _3625_ _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4534_ _1203_ _1098_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5137__C _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4465_ _0923_ _1135_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7253_ _3588_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _2771_ _2815_ _2818_ _2685_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7184_ _3547_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5510__A2 mod.Data_Mem.F_M.MRAM\[798\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4396_ _0647_ _0958_ _1063_ _1055_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _2186_ _2682_ _2750_ _1865_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_113_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6964__S _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ mod.Data_Mem.F_M.MRAM\[797\]\[0\] _2682_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5017_ _1681_ mod.Data_Mem.F_M.MRAM\[785\]\[1\] _1684_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7795__S _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6968_ _3405_ mod.Data_Mem.F_M.MRAM\[15\]\[7\] _3414_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5577__A2 mod.Data_Mem.F_M.MRAM\[799\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5919_ _1835_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6899_ mod.Data_Mem.F_M.dest\[4\] _3372_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6526__A1 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7574__I0 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6526__B2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8569_ _0073_ net349 mod.Data_Mem.F_M.out_data\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7326__I0 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8569__CLK net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6938__I _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__A2 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8077__D mod.P3.Res\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5265__A1 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6673__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5017__A1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4240__A2 mod.Arithmetic.CN.I_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8099__CLK net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8540__D _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6517__A1 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7565__I0 _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6517__B2 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ _0620_ _0922_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5343__I2 mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4181_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7940_ _0166_ net98 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6516__C _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7871_ _0097_ net372 mod.Data_Mem.F_M.MRAM\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5199__I _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6822_ mod.Data_Mem.F_M.MRAM\[789\]\[6\] _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _3283_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5927__I _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3965_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4862__S0 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5704_ _2065_ _2146_ _2329_ _2330_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_104_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6508__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6684_ _3228_ mod.Data_Mem.F_M.MRAM\[28\]\[0\] _3237_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8423_ _0519_ net92 mod.Data_Mem.F_M.MRAM\[790\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5635_ _2057_ _2111_ _2257_ _2267_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5863__S _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5031__I1 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8354_ _0450_ net292 mod.Data_Mem.F_M.MRAM\[781\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5566_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5731__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7305_ _3321_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4517_ mod.Arithmetic.CN.I_in\[12\] _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8285_ _0381_ net124 mod.Data_Mem.F_M.MRAM\[771\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5497_ _1835_ mod.Data_Mem.F_M.MRAM\[30\]\[5\] _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7236_ _3578_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4448_ _1111_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5495__A1 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7167_ _3538_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4379_ _0693_ _0810_ _1050_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6118_ _2732_ _2734_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7098_ mod.Data_Mem.F_M.MRAM\[23\]\[4\] _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6049_ _2635_ _2666_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5798__A2 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8241__CLK net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7795__I0 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4222__A2 mod.Arithmetic.CN.I_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4741__I _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8391__CLK net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7959__CLK net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A2 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5572__I _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5486__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5238__A1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4916__I _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6109__S _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__S1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7786__I0 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5261__I1 mod.Data_Mem.F_M.MRAM\[784\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout237_I net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__A2 mod.Data_Mem.F_M.MRAM\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6779__S _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _2076_ _0010_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5713__A2 mod.Data_Mem.F_M.MRAM\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5351_ _2008_ _2011_ _2013_ _1833_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4302_ _0952_ _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8070_ _0279_ net132 mod.Data_Mem.F_M.MRAM\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5282_ _1582_ _1945_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8114__CLK net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7021_ _3452_ mod.Data_Mem.F_M.MRAM\[18\]\[2\] _3448_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4233_ _0905_ _0906_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4164_ _0825_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_114_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4826__I mod.Data_Mem.F_M.src\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4095_ _0752_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8264__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7923_ _0149_ net122 mod.Data_Mem.F_M.MRAM\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4452__A2 mod.Arithmetic.CN.I_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7854_ _3929_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6805_ _3320_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7785_ _3890_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _1662_ _1663_ _1664_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6736_ _3273_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3948_ mod.P1.instr_reg\[17\] _0625_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6667_ mod.Data_Mem.F_M.MRAM\[27\]\[5\] _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8406_ _0502_ net97 mod.Data_Mem.F_M.MRAM\[787\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5618_ _2055_ mod.Data_Mem.F_M.MRAM\[797\]\[0\] _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5704__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ _3189_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6752__I1 mod.Data_Mem.F_M.MRAM\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8337_ _0433_ net211 mod.Data_Mem.F_M.MRAM\[778\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5392__I _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5549_ _2175_ _2182_ _2188_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8268_ _0364_ net127 mod.Data_Mem.F_M.MRAM\[768\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5468__A1 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7219_ _3568_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8199_ _0084_ net14 net114 mod.I_addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_48_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4140__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4443__A2 mod.Arithmetic.CN.I_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5640__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6951__I _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4672__S _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__A2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6172__B _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5567__I _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout60 net65 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout71 net72 net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5943__A2 mod.Data_Mem.F_M.MRAM\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3954__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout82 net83 net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout93 net94 net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6743__I1 mod.Data_Mem.F_M.MRAM\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8137__CLK net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4420__B _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4847__S _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6120__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7223__S _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout187_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7759__I0 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4851_ mod.Data_Mem.F_M.MRAM\[17\]\[0\] mod.Data_Mem.F_M.MRAM\[16\]\[0\] _1519_ _1520_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7570_ _3705_ _3335_ _3758_ _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4782_ _1447_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6521_ _2558_ mod.Data_Mem.F_M.MRAM\[780\]\[5\] _3115_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6452_ _2487_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5698__A1 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _2057_ _0010_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6383_ _2903_ mod.Data_Mem.F_M.MRAM\[15\]\[7\] mod.Data_Mem.F_M.MRAM\[14\]\[7\] _2253_
+ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8122_ mod.Data_Mem.F_M.out_data\[32\] net48 net337 mod.Arithmetic.CN.I_in\[32\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_126_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ _1888_ _1996_ _1624_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5145__C _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8053_ _0262_ net123 mod.Data_Mem.F_M.MRAM\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6111__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5265_ mod.Data_Mem.F_M.MRAM\[799\]\[4\] _1914_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7004_ _3441_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4216_ _0840_ _0889_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5196_ _1557_ _1825_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4147_ _0808_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4078_ _0681_ _0711_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__A2 mod.Arithmetic.CN.I_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5622__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5473__I1 mod.Data_Mem.F_M.MRAM\[799\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6771__I _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7906_ _0132_ net242 mod.Data_Mem.F_M.MRAM\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7837_ _3913_ _3915_ _3919_ _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_58_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7768_ _3880_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6719_ mod.Data_Mem.F_M.MRAM\[10\]\[2\] _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4984__I0 mod.Data_Mem.F_M.MRAM\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7699_ _3843_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5689__A1 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5689__B2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7107__I _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4361__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7043__S _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4113__A1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout250 net258 net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__B _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout261 net262 net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout272 net273 net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5861__A1 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout283 net284 net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout294 net295 net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8095__RN net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5613__A1 mod.Data_Mem.F_M.MRAM\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6681__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5613__B2 mod.Data_Mem.F_M.MRAM\[28\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5216__I1 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6964__I1 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7218__S _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7017__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout102_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7141__I1 mod.Data_Mem.F_M.MRAM\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5152__I0 mod.Data_Mem.F_M.MRAM\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _1610_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7841__A2 _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4001_ mod.P2.Rout_reg\[1\] _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5604__A1 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__B2 _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5952_ mod.Data_Mem.F_M.MRAM\[16\]\[5\] mod.Data_Mem.F_M.MRAM\[17\]\[5\] _2571_ _2572_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _1569_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5883_ _2338_ _1846_ _2504_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7622_ _3801_ _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4834_ mod.Data_Mem.F_M.src\[0\] _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5907__A2 mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout15_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7553_ _3759_ _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _1359_ _1360_ _1434_ _1358_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6032__S _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6504_ _3107_ _3108_ _2425_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7484_ _3292_ _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4696_ _1134_ _1251_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6435_ _2065_ _3041_ _3042_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6332__A2 _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5540__B1 mod.Data_Mem.F_M.MRAM\[798\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6366_ _2698_ _2023_ _2870_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8105_ mod.Data_Mem.F_M.out_data\[15\] net28 net268 mod.Arithmetic.CN.I_in\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4894__A2 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5317_ _1556_ _1980_ _1509_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7132__I1 mod.Data_Mem.F_M.MRAM\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6297_ mod.Data_Mem.F_M.MRAM\[781\]\[4\] _2745_ _2153_ mod.Data_Mem.F_M.MRAM\[780\]\[4\]
+ _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_88_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8036_ _0245_ net70 mod.Data_Mem.F_M.MRAM\[17\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5248_ _1557_ _1912_ _1863_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5843__A1 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5179_ _1514_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8077__RN net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7199__I1 mod.Data_Mem.F_M.MRAM\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6323__A2 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4334__A1 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__I _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5834__A1 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8325__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8543__D _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6562__A2 mod.Data_Mem.F_M.MRAM\[768\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout317_I net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4550_ _1122_ _1139_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__S _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6314__A2 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4481_ _1047_ _1084_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6220_ _1936_ _1818_ _2832_ _2833_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5373__I0 mod.Data_Mem.F_M.MRAM\[769\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _2708_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7114__I1 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _2698_ _1612_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ mod.Data_Mem.F_M.MRAM\[799\]\[1\] _1679_ _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4834__I mod.Data_Mem.F_M.src\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5589__B1 mod.Data_Mem.F_M.MRAM\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6984_ _3429_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5053__A2 mod.Data_Mem.F_M.MRAM\[769\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6250__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5935_ _1532_ _2135_ _2547_ _2554_ _2555_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _2487_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7050__I0 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7605_ _3754_ mod.Data_Mem.F_M.MRAM\[786\]\[5\] _3787_ _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0803_ _0678_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8585_ _0601_ net168 mod.Data_Mem.F_M.MRAM\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8231__RN net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6553__A2 mod.Data_Mem.F_M.MRAM\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ _2420_ mod.Data_Mem.F_M.MRAM\[789\]\[1\] _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7536_ _3711_ mod.Data_Mem.F_M.MRAM\[783\]\[3\] _3745_ _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4748_ _1414_ _1415_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7467_ _3708_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6305__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ _1225_ _1233_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7992__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6418_ _2346_ _2266_ _2358_ _3026_ _2354_ _2499_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7398_ _3672_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6349_ _1995_ _1994_ _1844_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6069__A1 mod.Data_Mem.F_M.MRAM\[781\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8019_ _0228_ net232 mod.Data_Mem.F_M.MRAM\[15\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5776__S _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7041__I0 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4555__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4307__B2 mod.Arithmetic.CN.I_in\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8538__D _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4919__I _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6480__A1 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__C _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7865__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3981_ _0649_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5720_ _2202_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4794__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__B1 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5651_ _2062_ _2282_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6535__A2 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4602_ _1149_ _1271_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4546__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8370_ _0466_ net292 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5582_ _1761_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7321_ _3630_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4533_ _1203_ _1099_ _1204_ _1095_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6299__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7252_ mod.Data_Mem.F_M.MRAM\[31\]\[2\] _3306_ _3585_ _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4464_ _0923_ _1019_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6203_ _2702_ _2816_ _2817_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7183_ mod.Data_Mem.F_M.MRAM\[22\]\[6\] _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4395_ _0956_ _1059_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _2744_ _2749_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _2674_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7141__S _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6471__A1 _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5016_ _1682_ _1683_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6980__S _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6223__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _3418_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5918_ _2259_ mod.Data_Mem.F_M.MRAM\[772\]\[4\] _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6898_ mod.Data_Mem.F_M.dest\[2\] _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5395__I _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5849_ _2425_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6526__A2 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8568_ _0072_ net340 mod.Data_Mem.F_M.out_data\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7519_ _3740_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7326__I1 mod.Data_Mem.F_M.MRAM\[770\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8499_ _0003_ net265 mod.Data_Mem.F_M.out_data\[75\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6837__I0 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7888__CLK net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6214__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4076__I0 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7785__I _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5973__B1 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7565__I1 mod.Data_Mem.F_M.MRAM\[784\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4528__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4700__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4180_ _0678_ _0679_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout384_I net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6453__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__B2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_560 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7870_ _0096_ net375 mod.Data_Mem.F_M.MRAM\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6205__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6821_ _3329_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _3259_ mod.Data_Mem.F_M.MRAM\[0\]\[7\] _3279_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4767__A1 mod.Arithmetic.CN.I_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3964_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7005__I0 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4862__S1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ _2169_ mod.Data_Mem.F_M.MRAM\[28\]\[6\] _2311_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6683_ _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_31_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8422_ _0518_ net86 mod.Data_Mem.F_M.MRAM\[790\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5148__C _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ _2067_ _2258_ _2266_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8353_ _0449_ net293 mod.Data_Mem.F_M.MRAM\[781\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5565_ _2202_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7304_ _3619_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4516_ _0621_ _0737_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8284_ _0380_ net110 mod.Data_Mem.F_M.MRAM\[771\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5496_ _1693_ mod.Data_Mem.F_M.MRAM\[798\]\[5\] _2139_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_89_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7235_ _3531_ mod.Data_Mem.F_M.MRAM\[30\]\[3\] _3574_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4447_ _1118_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5495__A2 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7166_ _3537_ mod.Data_Mem.F_M.MRAM\[12\]\[6\] _3534_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4378_ _0880_ _0954_ _0962_ _0963_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6117_ _1540_ _1516_ _1520_ _1614_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _3495_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ mod.Data_Mem.F_M.MRAM\[2\]\[7\] mod.Data_Mem.F_M.MRAM\[3\]\[7\] _2179_ _2666_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7244__I0 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7999_ _0208_ net305 mod.Data_Mem.F_M.MRAM\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7795__I1 mod.Data_Mem.F_M.MRAM\[798\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6442__C _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5183__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7046__S _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8088__D mod.P2.Rout_reg1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5486__A2 _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__A3 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5238__A2 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8066__CLK net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4997__A1 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7235__I0 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7786__I1 mod.Data_Mem.F_M.MRAM\[798\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4749__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__S _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout132_I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7903__CLK net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _1576_ _2012_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4301_ _0902_ _0970_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_114_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ mod.Data_Mem.F_M.MRAM\[787\]\[5\] mod.Data_Mem.F_M.MRAM\[786\]\[5\] _1944_
+ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6123__B1 mod.Data_Mem.F_M.MRAM\[782\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5316__I3 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _3242_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4232_ _0841_ _0850_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ _0833_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8409__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ _0754_ _0769_ _0770_ _0665_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7922_ _0148_ net125 mod.Data_Mem.F_M.MRAM\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5003__I _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7853_ mod.Data_Mem.F_M.MRAM\[9\]\[5\] _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout45_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8559__CLK net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6543__B _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6804_ mod.Data_Mem.F_M.MRAM\[799\]\[6\] _3319_ _3313_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4842__I _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7784_ _3293_ mod.Data_Mem.F_M.MRAM\[798\]\[0\] _3889_ _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4996_ _1564_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6735_ _3269_ _3270_ _3272_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3947_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6666_ _3223_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8405_ _0501_ net105 mod.Data_Mem.F_M.MRAM\[787\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5617_ _2220_ _2247_ _2250_ _2175_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6597_ mod.Data_Mem.F_M.MRAM\[11\]\[2\] _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6901__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8336_ _0432_ net155 mod.Data_Mem.F_M.MRAM\[778\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__C _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5548_ _1762_ _2187_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8267_ _0363_ net183 mod.Data_Mem.F_M.MRAM\[768\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5479_ _1806_ _2125_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5468__A2 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7218_ _3533_ mod.Data_Mem.F_M.MRAM\[2\]\[4\] _3567_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8198_ _0083_ net14 net118 mod.I_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5622__B _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7149_ _3526_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8089__CLK net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4752__I _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7926__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6172__C _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout50 net51 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout61 net62 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout72 net76 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout83 net84 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3954__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout94 net95 net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5156__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6353__B1 mod.Data_Mem.F_M.MRAM\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4903__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8546__D _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6408__A1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5092__B1 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7759__I1 mod.Data_Mem.F_M.MRAM\[796\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _1518_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout347_I net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _1174_ _1448_ _1449_ _1450_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ _2641_ mod.Data_Mem.F_M.MRAM\[781\]\[5\] _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _2100_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5698__A2 mod.Data_Mem.F_M.MRAM\[796\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5402_ _2062_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4103__S _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6382_ _2978_ _2981_ _2988_ _2991_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8121_ mod.Data_Mem.F_M.out_data\[31\] net40 net274 mod.Arithmetic.CN.I_in\[31\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5333_ _1992_ _1993_ _1994_ _1995_ _1896_ _1540_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_86_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8231__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8052_ _0261_ net123 mod.Data_Mem.F_M.MRAM\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ _1919_ _1928_ _1680_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7003_ _3399_ mod.Data_Mem.F_M.MRAM\[17\]\[4\] _3440_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4215_ _0829_ _0851_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _1624_ _1838_ _1860_ _1490_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4146_ _0816_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__S _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4077_ mod.Arithmetic.ACTI.x\[1\] _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7905_ _0131_ net307 mod.Data_Mem.F_M.MRAM\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7836_ _3907_ mod.I_addr\[2\] _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5386__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _1574_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7767_ _3303_ mod.Data_Mem.F_M.MRAM\[797\]\[1\] _3878_ _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6718_ _3262_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7698_ mod.Data_Mem.F_M.MRAM\[793\]\[1\] _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4984__I1 mod.Data_Mem.F_M.MRAM\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6649_ mod.Data_Mem.F_M.MRAM\[25\]\[4\] _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5689__A2 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8319_ _0415_ net79 mod.Data_Mem.F_M.MRAM\[775\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7324__S _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__B _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5352__B _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5310__A1 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout240 net241 net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout251 net253 net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout262 net285 net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout273 net283 net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout284 net285 net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout295 net326 net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5613__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6183__B _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__B1 mod.Data_Mem.F_M.MRAM\[782\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5301__A1 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5152__I1 mod.Data_Mem.F_M.MRAM\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6077__C _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4000_ _0653_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_65_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A2 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _1712_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4902_ mod.Data_Mem.F_M.MRAM\[773\]\[0\] mod.Data_Mem.F_M.MRAM\[772\]\[0\] _1570_
+ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5882_ _2503_ mod.Data_Mem.F_M.MRAM\[773\]\[3\] _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7601__I0 _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4833_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7621_ _3803_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7552_ _3761_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4764_ _1352_ _1361_ _1433_ _1226_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__C _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6503_ _2641_ mod.Data_Mem.F_M.MRAM\[769\]\[4\] _3058_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7483_ _3717_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4695_ mod.Arithmetic.CN.I_in\[62\] _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7208__I _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6434_ _2632_ mod.Data_Mem.F_M.MRAM\[13\]\[1\] _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5915__I0 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6365_ _2889_ _2022_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5540__A1 _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5540__B2 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5951__I _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8104_ mod.Data_Mem.F_M.out_data\[14\] net30 net269 mod.Arithmetic.CN.I_in\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5316_ _1976_ _1977_ _1978_ _1979_ _1526_ _1530_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6296_ _2746_ _2908_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7293__A1 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8035_ _0244_ net71 mod.Data_Mem.F_M.MRAM\[17\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6983__S _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _1905_ _1907_ _1909_ _1910_ _1911_ _1645_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6340__I0 mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5843__A2 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5178_ _1525_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4129_ _0665_ _0802_ _0804_ _0805_ _0628_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_56_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5151__S0 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8127__CLK net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7819_ mod.I_addr\[0\] mod.I_addr\[2\] mod.I_addr\[1\] _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4031__A1 mod.Arithmetic.CN.I_in\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4334__A2 mod.Arithmetic.CN.I_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5531__A1 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7054__S _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__A2 _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__A2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5302__S _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5598__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6011__A2 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4940__I _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5770__A1 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4573__A2 mod.Arithmetic.ACTI.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout212_I net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _1042_ _1150_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5373__I1 mod.Data_Mem.F_M.MRAM\[768\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5522__A1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5771__I _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5522__B2 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _1911_ _1668_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5101_ _1583_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _1588_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _1680_ _1699_ _1561_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__S _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5212__S _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5589__A1 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__S0 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6983_ _3399_ mod.Data_Mem.F_M.MRAM\[16\]\[4\] _3428_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5589__B2 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5011__I _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5934_ _2059_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__B1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5865_ _2388_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6551__B _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7139__S _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4850__I _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7604_ _3793_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7050__I1 mod.Data_Mem.F_M.MRAM\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4816_ _1395_ _1392_ _1484_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8584_ _0600_ net171 mod.Data_Mem.F_M.MRAM\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5796_ _1880_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6978__S _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _1373_ mod.Arithmetic.CN.I_in\[70\] _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5761__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7535_ _3750_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7466_ _3603_ mod.Data_Mem.F_M.MRAM\[780\]\[0\] _3707_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7990__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4678_ _1237_ _1256_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6417_ _2419_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7397_ mod.Data_Mem.F_M.MRAM\[774\]\[7\] _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6348_ _2867_ _2958_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6069__A2 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _2883_ _2886_ _2891_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6474__C1 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8018_ _0227_ net306 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4875__I0 mod.Data_Mem.F_M.MRAM\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5630__B _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7041__I1 mod.Data_Mem.F_M.MRAM\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__B1 mod.Data_Mem.F_M.MRAM\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4555__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6687__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5504__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4307__A2 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8554__D _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4491__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout162_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3980_ _0655_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4243__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8592__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__B2 _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5766__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _2277_ _2120_ _2279_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _1152_ _1260_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5581_ _2112_ _2213_ _2217_ _2218_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6791__I0 mod.Data_Mem.F_M.MRAM\[799\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7320_ _3615_ mod.Data_Mem.F_M.MRAM\[770\]\[4\] _3623_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4532_ _1101_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7251_ _3587_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4463_ _0616_ mod.Arithmetic.CN.I_in\[60\] _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _1733_ _1772_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ _3546_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4394_ _1058_ _1060_ _1065_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_98_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ mod.Data_Mem.F_M.MRAM\[13\]\[1\] _2745_ _2153_ mod.Data_Mem.F_M.MRAM\[12\]\[1\]
+ _2748_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5006__I _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout75_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _2170_ _2680_ _1731_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ mod.Data_Mem.F_M.MRAM\[784\]\[1\] _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4845__I _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6223__A2 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6966_ _3403_ mod.Data_Mem.F_M.MRAM\[15\]\[6\] _3414_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4234__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5917_ _2389_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4785__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6897_ _3334_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4580__I _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5609__C _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5848_ _2426_ _2466_ _2467_ _2431_ _2470_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4537__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8567_ _0071_ net247 mod.Data_Mem.F_M.out_data\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5779_ _2394_ _2403_ _2371_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7518_ _3725_ mod.Data_Mem.F_M.MRAM\[782\]\[4\] _3739_ _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8498_ _0002_ net339 mod.Data_Mem.F_M.out_data\[74\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7449_ mod.Data_Mem.F_M.MRAM\[778\]\[1\] _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5337__I1 mod.Data_Mem.F_M.MRAM\[768\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__I1 mod.Data_Mem.F_M.MRAM\[769\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8140__RN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6214__A2 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4776__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__B2 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4528__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6150__A1 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7242__S _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6366__B _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6453__A2 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8131__RN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout377_I net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_550 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_561 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6205__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6820_ mod.Data_Mem.F_M.MRAM\[789\]\[5\] _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7982__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6751_ _3282_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3963_ _0639_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ _2309_ mod.Data_Mem.F_M.MRAM\[29\]\[6\] _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6682_ _3230_ _3232_ _3235_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6359__I3 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8421_ _0517_ net162 mod.Data_Mem.F_M.MRAM\[790\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8198__RN net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ _2260_ _2263_ _2265_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4519__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__A1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5564_ _1553_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8352_ _0448_ net291 mod.Data_Mem.F_M.MRAM\[781\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5192__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7303_ _3618_ mod.Data_Mem.F_M.MRAM\[768\]\[6\] _3608_ _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4515_ _1166_ _1184_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8283_ _0379_ net296 mod.Data_Mem.F_M.MRAM\[771\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5495_ _1658_ mod.Data_Mem.F_M.MRAM\[799\]\[5\] _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7234_ _3577_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4446_ _0619_ _0930_ _0928_ _1114_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_132_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7165_ _3255_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4377_ _0962_ _0963_ _0879_ _0954_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_98_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _2700_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7096_ mod.Data_Mem.F_M.MRAM\[23\]\[3\] _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6047_ _2183_ _2150_ _2664_ _2258_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4455__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6790__I _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7244__I1 mod.Data_Mem.F_M.MRAM\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4207__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ mod.P2.dest_reg1\[8\] net25 net240 mod.P2.dest_reg\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5955__A1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__A2 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _3295_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5707__A1 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6132__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8113__RN net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7235__I1 mod.Data_Mem.F_M.MRAM\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5946__A1 _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4749__A2 mod.Arithmetic.CN.I_in\[70\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6994__I0 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6746__I0 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6371__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6371__B2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5265__B _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4300_ _0972_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5280_ _1583_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6123__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6123__B2 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4231_ _0841_ _0850_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5309__S0 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4162_ _0836_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__A1 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__A2 mod.Data_Mem.F_M.MRAM\[781\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8104__RN net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4093_ _0712_ _0757_ _0751_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__8010__CLK net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4437__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7921_ _0147_ net209 mod.Data_Mem.F_M.MRAM\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7852_ _3928_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6803_ _3318_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8160__CLK net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout38_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6985__I0 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7783_ _3888_ _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4995_ mod.Data_Mem.F_M.MRAM\[19\]\[1\] mod.Data_Mem.F_M.MRAM\[18\]\[1\] _1519_ _1663_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _3271_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3946_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6737__I0 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6665_ mod.Data_Mem.F_M.MRAM\[27\]\[4\] _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8404_ _0500_ net97 mod.Data_Mem.F_M.MRAM\[787\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5616_ mod.Data_Mem.F_M.MRAM\[797\]\[7\] _2221_ _2222_ mod.Data_Mem.F_M.MRAM\[796\]\[7\]
+ _2249_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_30_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6596_ _3188_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7878__CLK net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8335_ _0431_ net370 mod.Data_Mem.F_M.MRAM\[777\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5547_ _2165_ _2183_ _2155_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5890__S _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6114__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8266_ _0362_ net203 mod.Data_Mem.F_M.MRAM\[768\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5478_ _0025_ _2123_ _2124_ _2093_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6114__B2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6785__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7217_ _3561_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4429_ _1095_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8197_ _0082_ net15 net118 mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7148_ _3523_ mod.Data_Mem.F_M.MRAM\[12\]\[0\] _3525_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7079_ _3486_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4428__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__I0 mod.Data_Mem.F_M.MRAM\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8503__CLK net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5228__I0 mod.Data_Mem.F_M.MRAM\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6976__I0 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout40 net42 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout51 net68 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout62 net64 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout73 net75 net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout84 net94 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout95 net96 net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_80_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6353__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6353__B2 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4903__A2 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4116__B1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6695__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8033__CLK net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4667__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6408__A2 mod.Data_Mem.F_M.MRAM\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7520__S _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8562__D _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__B2 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4780_ _1310_ _1318_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4052__C1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6344__A1 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6450_ _2410_ _1775_ _3056_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5401_ _2061_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6381_ _2879_ _2989_ _2990_ _2897_ _1675_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ mod.Data_Mem.F_M.MRAM\[17\]\[6\] mod.Data_Mem.F_M.MRAM\[16\]\[6\] _1718_ _1995_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8120_ mod.Data_Mem.F_M.out_data\[30\] net41 net276 mod.Arithmetic.CN.I_in\[30\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8051_ _0260_ net125 mod.Data_Mem.F_M.MRAM\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5263_ _1920_ _1925_ _1927_ _1833_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4658__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7002_ _3434_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4214_ _0829_ _0851_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5194_ _1724_ _1850_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4145_ _0819_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5014__I _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__B1 mod.Data_Mem.F_M.MRAM\[798\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4076_ _0630_ _0710_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7904_ _0130_ net320 mod.Data_Mem.F_M.MRAM\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7835_ _3175_ _3918_ _3916_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6958__I0 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7766_ _3879_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4978_ mod.Data_Mem.F_M.MRAM\[6\]\[1\] _1643_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6717_ mod.Data_Mem.F_M.MRAM\[10\]\[1\] _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7697_ _3842_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6648_ _3214_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6335__A1 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6579_ _3177_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7605__S _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8318_ _0414_ net85 mod.Data_Mem.F_M.MRAM\[775\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7835__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8249_ _0345_ net314 mod.Data_Mem.F_M.MRAM\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout230 net231 net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5310__A2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout241 net260 net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout252 net253 net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout263 net285 net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout274 net276 net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout285 net286 net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout296 net300 net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__B _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7515__S _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4003__I mod.Arithmetic.CN.I_in\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8549__CLK net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8557__D _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4938__I _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout192_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7250__S _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5950_ _2447_ _2569_ _1536_ _2355_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_34_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4901_ _1543_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5881_ _1845_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7620_ _3765_ mod.Data_Mem.F_M.MRAM\[787\]\[3\] _3801_ _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4832_ mod.Data_Mem.F_M.src\[2\] _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6565__A1 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7551_ _3718_ mod.Data_Mem.F_M.MRAM\[784\]\[0\] _3760_ _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4763_ _1252_ _1354_ mod.Arithmetic.CN.I_in\[54\] _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8079__CLK net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _3084_ mod.Data_Mem.F_M.MRAM\[768\]\[4\] _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6317__A1 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7482_ _3620_ mod.Data_Mem.F_M.MRAM\[780\]\[7\] _3713_ _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4694_ _1250_ _1254_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ _2590_ mod.Data_Mem.F_M.MRAM\[12\]\[1\] _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5915__I1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7117__I0 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6364_ _2873_ _2020_ _2767_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5540__A2 mod.Data_Mem.F_M.MRAM\[799\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8103_ mod.Data_Mem.F_M.out_data\[13\] net30 net270 mod.Arithmetic.CN.I_in\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5315_ mod.Data_Mem.F_M.MRAM\[17\]\[5\] mod.Data_Mem.F_M.MRAM\[16\]\[5\] _1971_ _1979_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6295_ _2142_ mod.Data_Mem.F_M.MRAM\[783\]\[4\] mod.Data_Mem.F_M.MRAM\[782\]\[4\]
+ _1494_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8034_ _0243_ net210 mod.Data_Mem.F_M.MRAM\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7293__A2 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5246_ _1647_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5177_ _1839_ _1842_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4128_ _0801_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5679__I _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4103__I0 mod.Arithmetic.CN.I_in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4059_ _0685_ _0704_ _0719_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5151__S1 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4803__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7818_ mod.I_addr\[4\] mod.I_addr\[6\] mod.I_addr\[5\] mod.I_addr\[7\] _3908_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6556__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7749_ _3869_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4582__A3 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7108__I0 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5531__A2 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__B _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6973__I _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A1 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4022__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7309__I _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__I _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7347__I0 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8371__CLK net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5100_ _1704_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6080_ _2692_ _2694_ _2696_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__A1 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _1685_ _1688_ _1691_ _1697_ _1698_ _1565_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6982_ _3422_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5589__A2 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__S1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _2548_ _2549_ _2553_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6538__A1 _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5864_ _2484_ _2485_ _2371_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6538__B2 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7603_ _3778_ mod.Data_Mem.F_M.MRAM\[786\]\[4\] _3787_ _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout20_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4815_ _1395_ _1392_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8583_ _0599_ net101 mod.Instr_Mem.instruction\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5795_ _2388_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7534_ _3749_ mod.Data_Mem.F_M.MRAM\[783\]\[2\] _3745_ _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4746_ mod.Arithmetic.CN.I_in\[69\] _1376_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7465_ _3706_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5962__I _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4677_ _1238_ _1255_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6416_ _2535_ _3018_ _3024_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _3671_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6994__S _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6347_ _2954_ _2955_ _2956_ _2957_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _2713_ _2888_ _2890_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6474__B1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8017_ _0226_ net306 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6793__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6474__C2 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5229_ mod.Data_Mem.F_M.MRAM\[19\]\[4\] mod.Data_Mem.F_M.MRAM\[18\]\[4\] _1718_ _1894_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__I1 mod.Data_Mem.F_M.MRAM\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__B1 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8244__CLK net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5824__I0 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4252__A2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6529__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__B2 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8510__571 net571 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5504__A2 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5313__S _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8570__D _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout155_I net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6371__C _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__A2 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout322_I net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4600_ _1152_ _1260_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5580_ _2175_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5743__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6791__I1 _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6379__S0 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7250_ _1634_ _3303_ _3585_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4462_ _0661_ _1017_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8117__CLK net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6201_ _2774_ _1777_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7181_ mod.Data_Mem.F_M.MRAM\[22\]\[5\] _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4393_ _0633_ _0959_ _1062_ _1055_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_131_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _2746_ _2747_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6063_ _2679_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8267__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _1518_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout68_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5806__I0 mod.Data_Mem.F_M.MRAM\[782\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _3417_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5431__A1 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ mod.Data_Mem.F_M.MRAM\[770\]\[4\] mod.Data_Mem.F_M.MRAM\[771\]\[4\] _2490_
+ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7559__I0 _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6896_ _3370_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3993__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _2432_ _2468_ _2469_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6989__S _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8566_ _0070_ net248 mod.Data_Mem.F_M.out_data\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5778_ _2398_ _2402_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7517_ _3733_ _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4729_ _1280_ _1397_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8497_ _0001_ net268 mod.Data_Mem.F_M.out_data\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7448_ _3697_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7379_ mod.Data_Mem.F_M.MRAM\[773\]\[6\] _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7613__S _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4101__I _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4170__A1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3940__I _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4972__S _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5422__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6698__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5308__S _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5489__A1 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__I _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6150__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4011__I mod.Arithmetic.CN.I_in\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4161__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_540 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5978__S _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4464__A2 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_551 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5661__A1 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout272_I net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5413__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6750_ _3256_ mod.Data_Mem.F_M.MRAM\[0\]\[6\] _3279_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3962_ mod.Arithmetic.CN.F_in\[0\] _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output9_I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3975__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5701_ _2328_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _3234_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8420_ _0516_ net86 mod.Data_Mem.F_M.MRAM\[790\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5632_ _2264_ _2110_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4519__A3 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__A2 mod.Data_Mem.F_M.MRAM\[796\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8351_ _0447_ net229 mod.Data_Mem.F_M.MRAM\[780\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5563_ _2175_ _2192_ _2201_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7302_ _3318_ _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4514_ _1185_ _1093_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8282_ _0378_ net314 mod.Data_Mem.F_M.MRAM\[771\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5494_ _2118_ _2135_ _2138_ _2132_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7233_ _3529_ mod.Data_Mem.F_M.MRAM\[30\]\[2\] _3574_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4445_ _1112_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7164_ _3536_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4376_ _0966_ _0965_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6557__B _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6429__B1 _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4856__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ _2366_ _2684_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ _3494_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _2529_ _2657_ _2660_ _2663_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5652__A1 _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4455__A2 mod.Arithmetic.ACTI.x\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ mod.P2.dest_reg1\[4\] net20 net223 mod.P2.dest_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4207__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _3406_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5955__A2 _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6879_ mod.Data_Mem.F_M.MRAM\[6\]\[7\] _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5707__A2 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8549_ _0053_ net277 mod.Data_Mem.F_M.out_data\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3935__I mod.Arithmetic.CN.F_in\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4391__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4143__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4446__A2 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6994__I1 mod.Data_Mem.F_M.MRAM\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7518__S _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4006__I mod.Arithmetic.I_out\[79\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6746__I1 mod.Data_Mem.F_M.MRAM\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6371__A2 _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4382__A1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout118_I net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6123__A2 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4230_ _0843_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5882__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4161_ _0659_ mod.Arithmetic.CN.I_in\[40\] mod.Arithmetic.CN.I_in\[41\] _0837_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5309__S1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__A2 _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4092_ _0755_ _0768_ _0716_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5634__A1 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4437__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7920_ _0146_ net204 mod.Data_Mem.F_M.MRAM\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6891__I mod.Data_Mem.F_M.MRAM\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7851_ mod.Data_Mem.F_M.MRAM\[9\]\[4\] _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6802_ net9 _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7782_ _3294_ _3298_ _3446_ _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4994_ _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6985__I1 mod.Data_Mem.F_M.MRAM\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3948__A1 mod.P1.instr_reg\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6733_ mod.Data_Mem.F_M.dest\[4\] mod.Data_Mem.F_M.dest\[2\] _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3945_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4070__B1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _3222_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8455__CLK net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6737__I1 mod.Data_Mem.F_M.MRAM\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8403_ _0499_ net179 mod.Data_Mem.F_M.MRAM\[787\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5615_ _2223_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6595_ mod.Data_Mem.F_M.MRAM\[11\]\[1\] _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6362__A2 _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8334_ _0430_ net313 mod.Data_Mem.F_M.MRAM\[777\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5546_ mod.Data_Mem.F_M.MRAM\[29\]\[1\] _1539_ _1813_ mod.Data_Mem.F_M.MRAM\[28\]\[1\]
+ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_117_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8265_ _0361_ net203 mod.Data_Mem.F_M.MRAM\[768\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5970__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ mod.Data_Mem.F_M.MRAM\[798\]\[2\] mod.Data_Mem.F_M.MRAM\[799\]\[2\] _1892_
+ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7163__S _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7216_ _3566_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4428_ _1096_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8196_ _0081_ net14 net118 mod.I_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5873__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7147_ _3524_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4359_ _0787_ _0805_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7078_ mod.Data_Mem.F_M.MRAM\[21\]\[2\] _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5476__I1 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _2529_ _2644_ _2646_ _2426_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_86_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5228__I1 mod.Data_Mem.F_M.MRAM\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6976__I1 mod.Data_Mem.F_M.MRAM\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6050__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout30 net31 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout41 net42 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout52 net53 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout63 net65 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout74 net75 net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout85 net87 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout96 net137 net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6353__A2 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4116__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7972__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5813__C _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5864__A1 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__A1 mod.Data_Mem.F_M.MRAM\[797\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8098__RN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5616__B2 mod.Data_Mem.F_M.MRAM\[796\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5092__A2 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5120__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8478__CLK net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7248__S _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout235_I net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6344__A2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5400_ _2060_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6380_ _2045_ _2046_ _1804_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5331_ mod.Data_Mem.F_M.MRAM\[19\]\[6\] mod.Data_Mem.F_M.MRAM\[18\]\[6\] _1809_ _1994_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5790__I _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8050_ _0259_ net209 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5262_ _1576_ _1926_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7001_ _3439_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5855__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4658__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4213_ _0869_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5193_ _1808_ _1854_ _1858_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4144_ _0621_ mod.Arithmetic.CN.I_in\[8\] _0715_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_95_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__B2 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4075_ _0712_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_95_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout50_I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7903_ _0129_ net312 mod.Data_Mem.F_M.MRAM\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7834_ _0080_ _3171_ _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6958__I1 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7765_ _3293_ mod.Data_Mem.F_M.MRAM\[797\]\[0\] _3878_ _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4977_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6716_ _3261_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7696_ mod.Data_Mem.F_M.MRAM\[793\]\[0\] _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5218__S0 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6647_ mod.Data_Mem.F_M.MRAM\[25\]\[3\] _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4346__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7995__CLK net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6578_ _3175_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8317_ _0413_ net158 mod.Data_Mem.F_M.MRAM\[775\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5529_ _2168_ mod.Data_Mem.F_M.MRAM\[798\]\[0\] mod.Data_Mem.F_M.MRAM\[799\]\[0\]
+ _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6099__A1 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__I0 mod.Data_Mem.F_M.MRAM\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8248_ _0344_ net339 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5846__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8179_ _0289_ net206 mod.Data_Mem.F_M.MRAM\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout220 net222 net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout231 net232 net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout242 net243 net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout253 net257 net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout264 net267 net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7599__A1 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout275 net281 net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout286 net392 net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout297 net299 net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_19_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6271__A1 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__C1 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6326__A2 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4337__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5837__A1 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7531__S _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8573__D _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4954__I _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout185_I net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7868__CLK net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout352_I net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4900_ _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5880_ _2500_ _1851_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6014__A1 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _1496_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7550_ _3759_ _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4576__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _1410_ _1429_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_53_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ mod.Data_Mem.F_M.MRAM\[780\]\[4\] mod.Data_Mem.F_M.MRAM\[782\]\[4\] mod.Data_Mem.F_M.MRAM\[781\]\[4\]
+ _1902_ _2264_ _2338_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7481_ _3716_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6317__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ _1241_ _1249_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6432_ _2618_ _3031_ _3039_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6363_ _2887_ _2021_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7117__I1 mod.Data_Mem.F_M.MRAM\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5226__S _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8102_ mod.Data_Mem.F_M.out_data\[12\] net32 net247 mod.Arithmetic.CN.I_in\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5314_ mod.Data_Mem.F_M.MRAM\[19\]\[5\] mod.Data_Mem.F_M.MRAM\[18\]\[5\] _1604_ _1978_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6294_ mod.Data_Mem.F_M.MRAM\[13\]\[4\] _2900_ _2901_ mod.Data_Mem.F_M.MRAM\[12\]\[4\]
+ _2906_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_88_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5828__A1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8033_ _0242_ net301 mod.Data_Mem.F_M.MRAM\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5245_ mod.Data_Mem.F_M.MRAM\[771\]\[4\] mod.Data_Mem.F_M.MRAM\[770\]\[4\] _1831_
+ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4500__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5176_ _1840_ mod.Data_Mem.F_M.MRAM\[775\]\[3\] _1841_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4864__I mod.Data_Mem.F_M.src\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4127_ _0803_ _0753_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4103__I1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4058_ _0728_ _0727_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__S _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7817_ mod.I_addr\[3\] _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6556__A2 _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6800__I0 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8023__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4567__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7748_ _3747_ mod.Data_Mem.F_M.MRAM\[796\]\[1\] _3867_ _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7679_ _3833_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4104__I mod.Arithmetic.ACTI.x\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4319__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5367__I0 mod.Data_Mem.F_M.MRAM\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8173__CLK net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3943__I _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7108__I1 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7150__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6244__A1 _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A2 mod.Data_Mem.F_M.MRAM\[771\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8516__CLK net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7347__I1 mod.Data_Mem.F_M.MRAM\[771\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4014__I _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5358__I0 mod.Data_Mem.F_M.MRAM\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8568__D _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6180__B1 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout100_I net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7261__S _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__A2 _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ _1575_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__A1 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6981_ _3427_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4797__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5932_ _2550_ _2551_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_65_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ mod.Data_Mem.F_M.MRAM\[786\]\[3\] mod.Data_Mem.F_M.MRAM\[787\]\[3\] _2376_
+ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6538__A2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7602_ _3792_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4814_ _1396_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6404__I _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8582_ _0598_ net100 mod.Instr_Mem.instruction\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5794_ _2400_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8196__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout13_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7533_ _3305_ _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _0622_ mod.Arithmetic.CN.I_in\[71\] _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7464_ _3269_ _3705_ _3374_ _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4676_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5464__B _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6415_ _3020_ _2352_ _3021_ _3022_ _3023_ _2361_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7395_ mod.Data_Mem.F_M.MRAM\[774\]\[6\] _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6346_ _1920_ _1986_ _2733_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6277_ _2889_ _1909_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8016_ _0225_ net302 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5228_ mod.Data_Mem.F_M.MRAM\[21\]\[4\] mod.Data_Mem.F_M.MRAM\[20\]\[4\] _1892_ _1893_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6474__B2 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5159_ _1807_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6226__A1 _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__B2 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__A2 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5824__I1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4788__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8539__CLK net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3938__I _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A2 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4960__A1 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7145__I _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4009__I mod.Arithmetic.CN.I_in\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__B _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7906__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout315_I net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4530_ mod.Arithmetic.CN.I_in\[44\] _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6379__S1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ mod.Arithmetic.CN.I_in\[60\] _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6200_ _2772_ _1764_ _1765_ _1558_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4703__A1 mod.Arithmetic.CN.I_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7180_ _3545_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4392_ _1061_ _1063_ _1064_ _0873_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _2114_ mod.Data_Mem.F_M.MRAM\[14\]\[1\] mod.Data_Mem.F_M.MRAM\[15\]\[1\] _1944_
+ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_113_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A2 mod.Data_Mem.F_M.MRAM\[786\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _2678_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _1584_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5806__I1 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6964_ _3416_ mod.Data_Mem.F_M.MRAM\[15\]\[5\] _3414_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5431__A2 _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ mod.Data_Mem.F_M.MRAM\[782\]\[4\] _1902_ _2434_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6895_ mod.Data_Mem.F_M.MRAM\[4\]\[7\] _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5846_ _2434_ mod.Data_Mem.F_M.MRAM\[773\]\[2\] _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3993__A2 mod.Arithmetic.ACTI.x\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5195__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8565_ _0069_ net247 mod.Data_Mem.F_M.out_data\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5777_ _2399_ _2401_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7166__S _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7516_ _3738_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4728_ _1283_ _1387_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8496_ _0000_ net268 mod.Data_Mem.F_M.out_data\[72\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7447_ mod.Data_Mem.F_M.MRAM\[778\]\[0\] _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4659_ _1209_ _1207_ _1329_ _1218_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7378_ _3662_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ _2235_ _2238_ _2937_ _2940_ _2079_ _2784_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_88_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8211__CLK net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6447__A1 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4538__B _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__I _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__A2 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5088__C _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5186__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6383__B1 mod.Data_Mem.F_M.MRAM\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5489__A2 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5733__I0 mod.Data_Mem.F_M.MRAM\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4161__A2 mod.Arithmetic.CN.I_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5324__S _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6438__A1 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6438__B2 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A1 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_530 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_541 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7238__I0 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_552 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5661__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout265_I net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5413__A2 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3961_ _0636_ mod.Arithmetic.CN.I_in\[24\] _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5700_ _2077_ _2323_ _2327_ _2302_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ mod.Data_Mem.F_M.dest\[8\] _3233_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3975__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5631_ _2087_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5177__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8350_ _0446_ net229 mod.Data_Mem.F_M.MRAM\[780\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5562_ _1762_ _2200_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7301_ _3617_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4513_ _1090_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8281_ _0377_ net314 mod.Data_Mem.F_M.MRAM\[771\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5493_ _2136_ mod.Data_Mem.F_M.MRAM\[798\]\[4\] _2137_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8234__CLK net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7232_ _3576_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4444_ _0928_ _1113_ _1115_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7163_ _3508_ mod.Data_Mem.F_M.MRAM\[12\]\[5\] _3534_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4375_ _0968_ _0965_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6429__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6114_ _1506_ _1513_ _2730_ _1936_ _2727_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6429__B2 _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7094_ mod.Data_Mem.F_M.MRAM\[23\]\[2\] _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6129__I _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6045_ _2345_ _2662_ _2347_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7229__I0 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5652__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4872__I mod.Data_Mem.F_M.src\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7996_ mod.P2.dest_reg1\[2\] net20 net224 mod.P2.dest_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6947_ _3405_ mod.Data_Mem.F_M.MRAM\[14\]\[7\] _3400_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6878_ _3361_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5168__A1 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _2446_ _2452_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8548_ _0052_ net252 mod.Data_Mem.F_M.out_data\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6117__B1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4391__A2 mod.Arithmetic.CN.I_in\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8479_ _0575_ net238 mod.Data_Mem.F_M.MRAM\[797\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4143__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5144__S _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7468__I0 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5371__C _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__I _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A3 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__B1 mod.Data_Mem.F_M.MRAM\[782\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6108__B1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4382__A2 mod.Arithmetic.CN.I_in\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7534__S _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8576__D _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4160_ _0657_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5989__S _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout382_I net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4091_ _0765_ _0766_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__A2 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7850_ _3927_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _3317_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7781_ _3887_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _1580_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6732_ _3234_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3948__A2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3944_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4070__B2 mod.Arithmetic.CN.I_in\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6663_ mod.Data_Mem.F_M.MRAM\[27\]\[3\] _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4641__B _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7508__I _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5229__S _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ _2229_ mod.Data_Mem.F_M.MRAM\[799\]\[7\] mod.Data_Mem.F_M.MRAM\[798\]\[7\]
+ _2225_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8402_ _0498_ net182 mod.Data_Mem.F_M.MRAM\[787\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6594_ _3187_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8333_ _0429_ net308 mod.Data_Mem.F_M.MRAM\[777\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5570__A1 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5545_ _2008_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8264_ _0360_ net187 mod.Data_Mem.F_M.MRAM\[768\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5476_ mod.Data_Mem.F_M.MRAM\[30\]\[2\] mod.Data_Mem.F_M.MRAM\[31\]\[2\] _1682_ _2123_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5858__C1 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7215_ _3531_ mod.Data_Mem.F_M.MRAM\[2\]\[3\] _3562_ _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4427_ _1097_ _1098_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4867__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8195_ _0080_ net14 net118 mod.I_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6370__I0 _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7146_ _3269_ _3270_ _3374_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4358_ _0627_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7077_ _3485_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4289_ _0960_ _0961_ _0957_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _2378_ _2043_ _2645_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4816__B _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__B2 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7979_ _0205_ net89 mod.Data_Mem.F_M.MRAM\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4107__I _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout20 net22 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout31 net32 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout42 net45 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout53 net54 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout64 net65 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout75 net76 net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__3946__I _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout86 net87 net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_70_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout97 net99 net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4043__S _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7153__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6197__C _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5864__A2 _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7613__I0 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A2 mod.Data_Mem.F_M.MRAM\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4052__A1 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7328__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout130_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout228_I net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5552__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ mod.Data_Mem.F_M.MRAM\[21\]\[6\] mod.Data_Mem.F_M.MRAM\[20\]\[6\] _1892_ _1993_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ mod.Data_Mem.F_M.MRAM\[785\]\[4\] mod.Data_Mem.F_M.MRAM\[784\]\[4\] _1610_
+ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7000_ _3397_ mod.Data_Mem.F_M.MRAM\[17\]\[3\] _3435_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4212_ _0883_ _0886_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5192_ _1844_ _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4143_ _0631_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5607__A2 mod.Data_Mem.F_M.MRAM\[799\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4074_ _0741_ _0749_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_49_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7902_ _0128_ net307 mod.Data_Mem.F_M.MRAM\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6407__I _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7833_ _0081_ _3917_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7764_ _3877_ _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4976_ _1528_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ mod.Data_Mem.F_M.MRAM\[10\]\[0\] _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8572__CLK net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7695_ _3841_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5218__S1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6646_ _3213_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6577_ mod.I_addr\[0\] mod.I_addr\[2\] mod.I_addr\[1\] _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8316_ _0412_ net83 mod.Data_Mem.F_M.MRAM\[775\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5528_ _1711_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5146__I1 mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8247_ _0343_ net133 mod.Data_Mem.F_M.MRAM\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5846__A2 mod.Data_Mem.F_M.MRAM\[773\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout210 net211 net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_8178_ _0288_ net191 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout221 net222 net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout232 net234 net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout243 net244 net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_101_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7129_ _3514_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout254 net255 net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout265 net267 net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout276 net281 net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__7599__A2 _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout287 net289 net287 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout298 net299 net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5221__I _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4282__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__B1 _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__C2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7349__S _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__A1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__I0 mod.Data_Mem.F_M.MRAM\[784\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4337__A2 mod.Arithmetic.ACTI.x\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5837__A2 mod.Data_Mem.F_M.MRAM\[789\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5332__S _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout178_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8595__CLK net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7259__S _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6014__A2 mod.Data_Mem.F_M.MRAM\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4970__I _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout345_I net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4830_ _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4761_ _1286_ _1324_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5773__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6500_ _3096_ _2313_ _2603_ _2546_ _3104_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7480_ _3618_ mod.Data_Mem.F_M.MRAM\[780\]\[6\] _3713_ _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _1350_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6431_ _2693_ _3038_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _2864_ _2972_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8101_ mod.Data_Mem.F_M.out_data\[11\] net36 net282 mod.Arithmetic.CN.I_in\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5313_ mod.Data_Mem.F_M.MRAM\[21\]\[5\] mod.Data_Mem.F_M.MRAM\[20\]\[5\] _1570_ _1977_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6293_ _2902_ _2905_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8032_ _0241_ net211 mod.Data_Mem.F_M.MRAM\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5244_ mod.Data_Mem.F_M.MRAM\[769\]\[4\] mod.Data_Mem.F_M.MRAM\[768\]\[4\] _1908_
+ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6340__I3 mod.Data_Mem.F_M.MRAM\[788\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _1704_ mod.Data_Mem.F_M.MRAM\[774\]\[3\] _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4500__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5242__S _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4126_ mod.P2.Rout_reg\[0\] _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6137__I _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4057_ _0731_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7169__S _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6005__A2 mod.Data_Mem.F_M.MRAM\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7816_ _3906_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6800__I1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__A2 mod.Arithmetic.CN.I_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7747_ _3868_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _1627_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7993__RN net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7678_ mod.Data_Mem.F_M.MRAM\[791\]\[7\] _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6629_ mod.Data_Mem.F_M.MRAM\[26\]\[2\] _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5367__I1 mod.Data_Mem.F_M.MRAM\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5660__B _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5152__S _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4991__S _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7744__A2 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5755__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4558__A2 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5507__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5358__I1 mod.Data_Mem.F_M.MRAM\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6180__A1 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6180__B2 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7542__S _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__I _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8161__RN net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6483__A2 mod.Data_Mem.F_M.MRAM\[780\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout295_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4494__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__C _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6980_ _3397_ mod.Data_Mem.F_M.MRAM\[16\]\[3\] _3423_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7985__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5931_ _2269_ mod.Data_Mem.F_M.MRAM\[20\]\[4\] _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4797__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5994__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5796__I _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5862_ _2381_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__I3 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7601_ _3765_ mod.Data_Mem.F_M.MRAM\[786\]\[3\] _3787_ _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4813_ _1399_ _1474_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8581_ _0597_ net218 mod.Instr_Mem.instruction\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5793_ _2296_ _1683_ _2416_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4205__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7532_ _3748_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4744_ _0622_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7463_ _3297_ _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5349__I1 mod.Data_Mem.F_M.MRAM\[784\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4675_ _1330_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6414_ _2487_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6171__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7394_ _3670_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6345_ _2873_ _1985_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5036__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6276_ _1581_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8015_ _0224_ net303 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5227_ _1610_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__6474__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _1808_ _1811_ _1814_ _1823_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_111_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109_ _0731_ _0784_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_5089_ _1509_ _1743_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5985__A1 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4788__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5737__A1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4115__I mod.Arithmetic.ACTI.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4960__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__A1 _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6486__B _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6465__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5976__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4453__C mod.Arithmetic.ACTI.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4400__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4951__A2 _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7336__I _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout210_I net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6240__I mod.Data_Mem.F_M.MRAM\[781\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout308_I net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4460_ _1124_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6153__A1 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4391_ _0613_ mod.Arithmetic.CN.I_in\[27\] _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6130_ _1525_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8134__RN net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6061_ _1710_ _2368_ _1496_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _1597_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6208__A2 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6963_ _3252_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8163__CLK net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5967__A1 _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _2098_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6894_ _3369_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5845_ _2209_ mod.Data_Mem.F_M.MRAM\[772\]\[2\] _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8564_ _0068_ net248 mod.Data_Mem.F_M.out_data\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5776_ mod.Data_Mem.F_M.MRAM\[786\]\[0\] mod.Data_Mem.F_M.MRAM\[787\]\[0\] _2400_
+ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7515_ _3711_ mod.Data_Mem.F_M.MRAM\[782\]\[3\] _3734_ _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4727_ _1283_ _1387_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8495_ _0591_ net72 mod.Data_Mem.F_M.MRAM\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7446_ _3696_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4658_ _1206_ _1213_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7377_ mod.Data_Mem.F_M.MRAM\[773\]\[5\] _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _1149_ _1152_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_89_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ mod.Data_Mem.F_M.MRAM\[781\]\[5\] _2745_ _2153_ mod.Data_Mem.F_M.MRAM\[780\]\[5\]
+ _2939_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5922__C _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8125__RN net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6447__A2 mod.Data_Mem.F_M.MRAM\[781\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6259_ _2855_ _1881_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4458__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4538__C _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__A1 _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6383__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5186__A2 _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6383__B2 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7156__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5733__I1 mod.Data_Mem.F_M.MRAM\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8036__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4161__A3 mod.Arithmetic.CN.I_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6438__A2 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8116__RN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4449__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A2 mod.Data_Mem.F_M.MRAM\[769\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_520 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_531 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_542 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7238__I1 mod.Data_Mem.F_M.MRAM\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_553 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5340__S _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout160_I net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5413__A3 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout258_I net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3960_ mod.Arithmetic.CN.I_in\[16\] _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4621__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5630_ _2261_ mod.Data_Mem.F_M.MRAM\[28\]\[0\] _2262_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8517__568 net568 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6374__A1 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5561_ _2155_ _2199_ _1632_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7066__I mod.Data_Mem.F_M.MRAM\[20\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7300_ _3569_ mod.Data_Mem.F_M.MRAM\[768\]\[5\] _3608_ _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4512_ _1169_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8280_ _0376_ net296 mod.Data_Mem.F_M.MRAM\[771\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5492_ _1615_ mod.Data_Mem.F_M.MRAM\[799\]\[4\] _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7231_ _3527_ mod.Data_Mem.F_M.MRAM\[30\]\[1\] _3574_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6677__A2 mod.Data_Mem.F_M.dest\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ _0632_ mod.Arithmetic.CN.I_in\[52\] _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5885__B1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7162_ _3535_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4374_ _0970_ _0974_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6113_ mod.Data_Mem.F_M.MRAM\[23\]\[0\] mod.Data_Mem.F_M.MRAM\[22\]\[0\] _1717_ _2730_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8107__RN net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7093_ _3493_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _2278_ mod.Data_Mem.F_M.MRAM\[18\]\[7\] _2661_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5732__S0 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7229__I1 mod.Data_Mem.F_M.MRAM\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7995_ mod.P2.dest_reg1\[1\] net19 net226 mod.P2.dest_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _3258_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6877_ mod.Data_Mem.F_M.MRAM\[6\]\[6\] _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5984__I _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6365__A1 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5168__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5828_ _2447_ _2451_ _1807_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8547_ _0051_ net327 mod.Data_Mem.F_M.out_data\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5759_ _2381_ _2382_ _2383_ _2273_ _2369_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8059__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6117__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8478_ _0574_ net237 mod.Data_Mem.F_M.MRAM\[797\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6117__B2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7429_ mod.Data_Mem.F_M.MRAM\[776\]\[7\] _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6912__I0 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7468__I1 mod.Data_Mem.F_M.MRAM\[780\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5224__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4446__A4 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5160__S _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A4 _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__I _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6108__A1 mod.Data_Mem.F_M.MRAM\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6108__B2 mod.Data_Mem.F_M.MRAM\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4119__B1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__B _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6903__I0 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _0750_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6292__B1 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout375_I net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5634__A3 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5890__I0 mod.Data_Mem.F_M.MRAM\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_394 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6800_ mod.Data_Mem.F_M.MRAM\[799\]\[5\] _3316_ _3313_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7780_ _3784_ mod.Data_Mem.F_M.MRAM\[797\]\[7\] _3883_ _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5398__A2 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ _1657_ _1659_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6731_ _3231_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3943_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6662_ _3221_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8201__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8401_ _0497_ net182 mod.Data_Mem.F_M.MRAM\[787\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ mod.Data_Mem.F_M.MRAM\[29\]\[7\] _2082_ _1642_ mod.Data_Mem.F_M.MRAM\[28\]\[7\]
+ _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ mod.Data_Mem.F_M.MRAM\[11\]\[0\] _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8332_ _0428_ net210 mod.Data_Mem.F_M.MRAM\[777\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5544_ _2088_ mod.Data_Mem.F_M.MRAM\[30\]\[1\] _1634_ _1954_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5570__A2 mod.Data_Mem.F_M.MRAM\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8263_ _0359_ net82 mod.Data_Mem.F_M.MRAM\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5475_ _2068_ _2117_ _2118_ _2120_ _2122_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5245__S _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5858__B1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7214_ _3565_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5858__C2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4426_ _0837_ _1097_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8194_ net574 net47 net333 mod.Arithmetic.CN.F_in\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_67_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7145_ _3227_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4357_ _0629_ _1028_ _1030_ mod.P3.Res\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4288_ _0957_ _0960_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_7076_ mod.Data_Mem.F_M.MRAM\[21\]\[1\] _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4883__I mod.Data_Mem.F_M.src\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6027_ _2196_ mod.Data_Mem.F_M.MRAM\[786\]\[7\] _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7978_ _0204_ net81 mod.Data_Mem.F_M.MRAM\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _3393_ mod.Data_Mem.F_M.MRAM\[14\]\[1\] _3391_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout21 net22 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout32 net33 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout43 net45 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6338__A1 _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout54 net67 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout65 net66 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout76 net77 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout87 net90 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout98 net99 net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5219__I _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3962__I mod.Arithmetic.CN.F_in\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6510__A1 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7310__I0 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6494__B _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5838__B _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4052__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8374__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5129__I _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5001__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout123_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5573__B _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5260_ _1921_ _1922_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4211_ mod.Arithmetic.CN.I_in\[8\] _0713_ _0818_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5191_ _1845_ mod.Data_Mem.F_M.MRAM\[769\]\[3\] _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4142_ _0817_ _0715_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4073_ mod.Arithmetic.CN.I_in\[15\] _0711_ _0747_ _0744_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_83_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7901_ _0127_ net303 mod.Data_Mem.F_M.MRAM\[27\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7832_ _3916_ _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout36_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7763_ _3230_ _3705_ _3371_ _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4975_ _1642_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6714_ _3260_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7694_ mod.Data_Mem.F_M.MRAM\[792\]\[7\] _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6645_ mod.Data_Mem.F_M.MRAM\[25\]\[2\] _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ _3174_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4346__A3 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8315_ _0411_ net142 mod.Data_Mem.F_M.MRAM\[775\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8246_ _0342_ net133 mod.Data_Mem.F_M.MRAM\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7296__A2 _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5458_ _2063_ _2058_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout200 net214 net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4409_ _1078_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8177_ mod.P1.instr_reg\[8\] net34 net261 mod.P2.Rout_reg1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout211 net212 net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5389_ _2034_ _2040_ _2050_ _1931_ _1630_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout222 net228 net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout233 net234 net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7128_ _3445_ mod.Data_Mem.F_M.MRAM\[19\]\[0\] _3513_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout244 net250 net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout255 net257 net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout266 net267 net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout277 net280 net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout288 net290 net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout299 net300 net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7059_ _3476_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4282__A2 mod.Arithmetic.CN.I_in\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A1 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6559__B2 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4034__A2 mod.Arithmetic.I_out\[79\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3957__I _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5909__I1 mod.Data_Mem.F_M.MRAM\[785\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6031__I0 mod.Data_Mem.F_M.MRAM\[782\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7531__I0 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5298__A1 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6709__S _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5412__I _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5222__A1 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout240_I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout338_I net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4760_ _1287_ _1323_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6970__A1 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5773__A2 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _1352_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _1536_ _3032_ _3034_ _3037_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6361_ _2866_ _2963_ _2971_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8100_ mod.Data_Mem.F_M.out_data\[10\] net58 net345 mod.Arithmetic.CN.I_in\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5312_ mod.Data_Mem.F_M.MRAM\[23\]\[5\] mod.Data_Mem.F_M.MRAM\[22\]\[5\] _1971_ _1976_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7522__I0 _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6292_ _2903_ mod.Data_Mem.F_M.MRAM\[15\]\[4\] mod.Data_Mem.F_M.MRAM\[14\]\[4\] _2904_
+ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8031_ _0240_ net210 mod.Data_Mem.F_M.MRAM\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5243_ _1514_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5174_ _1692_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4125_ _0678_ _0679_ _0801_ mod.P2.Rout_reg\[0\] _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_56_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4056_ _0732_ _0696_ _0719_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7815_ mod.Data_Mem.F_M.MRAM\[7\]\[7\] _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7746_ _3771_ mod.Data_Mem.F_M.MRAM\[796\]\[0\] _3867_ _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4958_ _1502_ _1533_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5992__I _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7677_ _3832_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4889_ _1552_ _1537_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6628_ _3204_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4319__A3 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__I0 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6559_ _3030_ _2343_ _3023_ _2646_ _2644_ _2484_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_106_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8229_ mod.P1.instr_reg\[11\] net17 net224 mod.P2.dest_reg1\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6264__S _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__B _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5204__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__I _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6004__I0 mod.Data_Mem.F_M.MRAM\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A2 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7752__I0 _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__I _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6180__A2 mod.Data_Mem.F_M.MRAM\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7622__I _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5691__A1 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4494__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout190_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8562__CLK net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5818__I0 mod.Data_Mem.F_M.MRAM\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4981__I _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5930_ _2304_ mod.Data_Mem.F_M.MRAM\[21\]\[4\] _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5994__A2 mod.Data_Mem.F_M.MRAM\[782\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _2081_ _2473_ _2483_ _1499_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7600_ _1793_ _3789_ _3791_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4812_ _1477_ _1479_ _1481_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8580_ _0596_ net119 mod.Instr_Mem.instruction\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5792_ _2075_ mod.Data_Mem.F_M.MRAM\[785\]\[1\] _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7531_ _3747_ mod.Data_Mem.F_M.MRAM\[783\]\[1\] _3745_ _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4743_ mod.Arithmetic.CN.I_in\[47\] _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7462_ _3704_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4674_ _1235_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6413_ _2381_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7393_ mod.Data_Mem.F_M.MRAM\[774\]\[5\] _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6171__A2 _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4182__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6344_ _1662_ _1987_ _2782_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6349__S _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6275_ _2887_ _1910_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8014_ _0223_ net126 mod.Data_Mem.F_M.MRAM\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5226_ mod.Data_Mem.F_M.MRAM\[23\]\[4\] mod.Data_Mem.F_M.MRAM\[22\]\[4\] _1890_ _1891_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4377__B _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4485__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ _1655_ _1817_ _1822_ _1645_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ _0733_ _0772_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5088_ _1745_ _1749_ _1751_ _1754_ _1619_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5434__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5985__A2 mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3996__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5737__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7729_ _3858_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4173__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3970__I _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5673__A1 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6058__I _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5976__A2 mod.Data_Mem.F_M.MRAM\[789\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__I _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5338__S _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4400__A2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout203_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4390_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4976__I _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _2675_ _2676_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ _1678_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6962_ _3415_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5913_ _2524_ _2138_ _2525_ _2528_ _2533_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6893_ mod.Data_Mem.F_M.MRAM\[4\]\[6\] _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ mod.Data_Mem.F_M.MRAM\[782\]\[2\] mod.Data_Mem.F_M.MRAM\[783\]\[2\] _1954_
+ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8563_ _0067_ net337 mod.Data_Mem.F_M.out_data\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ _1584_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6392__A2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7527__I _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7514_ _3737_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4726_ _1277_ _1388_ _1389_ _1274_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8494_ _0590_ net80 mod.Data_Mem.F_M.MRAM\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7445_ mod.Data_Mem.F_M.MRAM\[777\]\[7\] _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4657_ _1220_ _1326_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7376_ _3661_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4588_ _1154_ _1158_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_116_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6327_ _2746_ _2938_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6258_ _2698_ _1877_ _2870_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5655__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _1873_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _2178_ _1738_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6383__A2 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3965__I _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6135__A2 _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4146__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6497__B _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4449__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_510 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_521 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_532 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_543 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_554 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4036__I mod.Arithmetic.CN.I_in\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout153_I net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout320_I net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6251__I _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ mod.Data_Mem.F_M.MRAM\[29\]\[2\] _2193_ _2195_ mod.Data_Mem.F_M.MRAM\[28\]\[2\]
+ _2198_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4511_ _1058_ _1172_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5491_ _1692_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6126__A2 _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7230_ _3575_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4442_ mod.Arithmetic.CN.I_in\[50\] _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5885__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7161_ _3533_ mod.Data_Mem.F_M.MRAM\[12\]\[4\] _3534_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5885__B2 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7082__I mod.Data_Mem.F_M.MRAM\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4373_ _1044_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6112_ _2366_ _2680_ _2724_ _2725_ _2728_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_112_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7092_ mod.Data_Mem.F_M.MRAM\[23\]\[1\] _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8130__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _1792_ mod.Data_Mem.F_M.MRAM\[19\]\[7\] _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5732__S1 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout66_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6437__I0 mod.Data_Mem.F_M.MRAM\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7994_ mod.P2.dest_reg1\[0\] net17 net223 mod.P2.dest_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _3404_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4073__B1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _3360_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5827_ _2448_ _2444_ _2350_ _2449_ _2450_ _2168_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4376__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7998__CLK net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8546_ _0050_ net331 mod.Data_Mem.F_M.out_data\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5758_ mod.Data_Mem.F_M.MRAM\[772\]\[0\] mod.Data_Mem.F_M.MRAM\[773\]\[0\] _1515_
+ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _1373_ _1379_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7314__A1 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8477_ _0573_ net235 mod.Data_Mem.F_M.MRAM\[797\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6117__A2 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ _2077_ _2313_ _2317_ _2302_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_159_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7428_ _3687_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7359_ mod.Data_Mem.F_M.MRAM\[772\]\[4\] _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A1 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4603__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6356__A2 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8003__CLK net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6108__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4119__B2 mod.Arithmetic.ACTI.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6903__I1 mod.Data_Mem.F_M.MRAM\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8153__CLK net361 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5415__I _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6292__A1 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5890__I1 mod.Data_Mem.F_M.MRAM\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout270_I net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout368_I net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_395 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6044__A1 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ mod.Data_Mem.F_M.MRAM\[17\]\[1\] mod.Data_Mem.F_M.MRAM\[16\]\[1\] _1658_ _1659_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6730_ _3268_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3942_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_output7_I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6661_ mod.Data_Mem.F_M.MRAM\[27\]\[2\] _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5612_ _1661_ _2245_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8400_ _0496_ net179 mod.Data_Mem.F_M.MRAM\[787\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6592_ _3186_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8331_ _0427_ net172 mod.Data_Mem.F_M.MRAM\[777\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ _1532_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8262_ _0358_ net91 mod.Data_Mem.F_M.MRAM\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5474_ _2093_ _2121_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5858__A1 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7213_ _3529_ mod.Data_Mem.F_M.MRAM\[2\]\[2\] _3562_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4425_ _0834_ mod.Arithmetic.CN.I_in\[41\] _0898_ _0984_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5858__B2 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8193_ _0303_ net109 mod.Data_Mem.F_M.MRAM\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7144_ _3522_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4356_ _0781_ _0857_ _0858_ _1029_ _0627_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_98_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7075_ _3484_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4287_ _0648_ _0959_ _0812_ _0875_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_98_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6026_ mod.Data_Mem.F_M.MRAM\[784\]\[7\] mod.Data_Mem.F_M.MRAM\[785\]\[7\] _2297_
+ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5330__I0 mod.Data_Mem.F_M.MRAM\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6156__I _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5060__I _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7977_ _0203_ net184 mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _3239_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout11 net13 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout22 net23 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout33 net37 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout44 net50 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6859_ mod.Data_Mem.F_M.MRAM\[779\]\[5\] _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout55 net56 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout66 net67 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout77 net96 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4349__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout88 net89 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5546__B1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout99 net103 net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8176__CLK net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8529_ _0033_ net332 mod.Data_Mem.F_M.out_data\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5849__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6510__A2 mod.Data_Mem.F_M.MRAM\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6267__S _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__A2 mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8519__CLK net361 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7526__A1 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5001__A2 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout116_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7561__S _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4210_ mod.Arithmetic.CN.I_in\[8\] _0818_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4512__A1 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5190_ _1649_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4141_ _0636_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5081__S _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4072_ _0742_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_77_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7900_ _0126_ net172 mod.Data_Mem.F_M.MRAM\[27\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7831_ _0612_ _3175_ _3916_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4028__B1 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6704__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7762_ _3876_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4974_ _1599_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8199__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6713_ _3259_ mod.Data_Mem.F_M.MRAM\[28\]\[7\] _3250_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7693_ _3840_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout29_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6644_ _3212_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5379__I0 mod.Data_Mem.F_M.MRAM\[791\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6575_ mod.I_addr\[3\] _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8314_ _0410_ net191 mod.Data_Mem.F_M.MRAM\[775\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5526_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8245_ _0341_ net132 mod.Data_Mem.F_M.MRAM\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5457_ _2105_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4408_ _0722_ _0820_ _0972_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8176_ mod.P1.instr_reg\[7\] net38 net262 mod.P2.Rout_reg1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5700__B1 _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout201 net202 net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_5388_ mod.Data_Mem.F_M.MRAM\[799\]\[7\] _1914_ _2049_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout212 net213 net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout223 net225 net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_7127_ _3512_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout234 net241 net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4339_ _1010_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout245 net249 net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout256 net257 net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout267 net272 net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6256__A1 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout278 net280 net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7058_ mod.Data_Mem.F_M.MRAM\[20\]\[0\] _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout289 net290 net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _2055_ mod.Data_Mem.F_M.MRAM\[18\]\[6\] _2627_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5004__B _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6008__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7056__I0 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A2 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4134__I _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6031__I1 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5166__S _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4742__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6495__A1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7531__I1 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7039__A3 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5222__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4044__I mod.Arithmetic.CN.I_in\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout233_I net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8491__CLK net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4690_ _1359_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4979__I _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4033__I0 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6360_ _2865_ _2970_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4733__A1 mod.Arithmetic.CN.I_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ mod.Data_Mem.F_M.MRAM\[31\]\[5\] _1934_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6291_ _1493_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7522__I1 mod.Data_Mem.F_M.MRAM\[782\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8030_ _0239_ net73 mod.Data_Mem.F_M.MRAM\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6486__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ mod.Data_Mem.F_M.MRAM\[775\]\[4\] mod.Data_Mem.F_M.MRAM\[774\]\[4\] _1906_
+ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5173_ _1647_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_96_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4124_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4219__I mod.Arithmetic.CN.I_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 io_in[8] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4055_ _0697_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5997__B1 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4663__B _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7814_ _3905_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7745_ _3866_ _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4957_ _1621_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7466__S _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6370__S _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7676_ mod.Data_Mem.F_M.MRAM\[791\]\[6\] _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4888_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6627_ mod.Data_Mem.F_M.MRAM\[26\]\[1\] _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6174__B1 mod.Data_Mem.F_M.MRAM\[782\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7265__I mod.Data_Mem.F_M.MRAM\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7761__I1 mod.Data_Mem.F_M.MRAM\[796\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4724__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _3096_ _2340_ _2657_ _3063_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ _1809_ mod.Data_Mem.F_M.MRAM\[799\]\[7\] _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6489_ _3083_ _3092_ _3094_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7513__I1 mod.Data_Mem.F_M.MRAM\[782\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8228_ mod.P1.instr_reg\[10\] net19 net219 mod.P2.dest_reg1\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8159_ mod.Data_Mem.F_M.out_data\[69\] net62 net358 mod.Arithmetic.CN.I_in\[69\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5513__I _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6229__A1 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5204__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6401__A1 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7201__I0 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6004__I1 mod.Data_Mem.F_M.MRAM\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7175__I mod.Data_Mem.F_M.MRAM\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5912__B1 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6012__C _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4191__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6468__A1 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5423__I _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5691__A2 mod.Data_Mem.F_M.MRAM\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5818__I1 mod.Data_Mem.F_M.MRAM\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4039__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout183_I net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5979__B1 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__A2 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout350_I net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6254__I _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5860_ _2478_ _2482_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _1363_ _1383_ _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7530_ _3302_ _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4742_ _1411_ mod.Arithmetic.CN.I_in\[46\] _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7461_ mod.Data_Mem.F_M.MRAM\[778\]\[7\] _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4673_ _1335_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6412_ mod.Data_Mem.F_M.MRAM\[0\]\[0\] mod.Data_Mem.F_M.MRAM\[1\]\[0\] _2705_ _3021_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8237__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4706__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7392_ _3669_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6343_ _2855_ _1988_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6459__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6274_ _1637_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout96_I net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8013_ _0222_ net126 mod.Data_Mem.F_M.MRAM\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5225_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5131__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7259__I0 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5156_ _1560_ _1819_ _1821_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4107_ _0752_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ _1752_ _1753_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ mod.Arithmetic.CN.I_in\[9\] _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3996__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5817__S0 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5198__A1 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ mod.Data_Mem.F_M.MRAM\[784\]\[6\] mod.Data_Mem.F_M.MRAM\[785\]\[6\] _2297_
+ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7728_ mod.Data_Mem.F_M.MRAM\[795\]\[0\] _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7659_ _3823_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5370__A1 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4173__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5122__A1 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5673__A2 mod.Data_Mem.F_M.MRAM\[797\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6386__B1 mod.Data_Mem.F_M.MRAM\[782\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6802__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6138__B1 mod.Data_Mem.F_M.MRAM\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__I0 mod.Data_Mem.F_M.MRAM\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5897__C1 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7489__I0 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _1596_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5664__A2 _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6961_ _3399_ _1870_ _3414_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__C1 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5912_ _2529_ _2530_ _2532_ _2426_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_35_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6892_ _3368_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ _2464_ _1770_ _2465_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8562_ _0066_ net347 mod.Data_Mem.F_M.out_data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5774_ _2107_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout11_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7513_ _3640_ mod.Data_Mem.F_M.MRAM\[782\]\[2\] _3734_ _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4725_ _1273_ _1390_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8493_ _0589_ net160 mod.Data_Mem.F_M.MRAM\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7444_ _3695_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4656_ _1223_ _1257_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5727__I0 mod.Data_Mem.F_M.MRAM\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4155__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7375_ mod.Data_Mem.F_M.MRAM\[773\]\[4\] _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4587_ _1197_ _1201_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6326_ _2268_ mod.Data_Mem.F_M.MRAM\[783\]\[5\] mod.Data_Mem.F_M.MRAM\[782\]\[5\]
+ _2904_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5104__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6257_ _2700_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5063__I _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5655__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5208_ _1583_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6188_ _1752_ _1741_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5998__I _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5139_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4918__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A1 mod.Data_Mem.F_M.MRAM\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4394__A2 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5591__B2 mod.Data_Mem.F_M.MRAM\[28\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3981__I _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6497__C _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_500 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_94_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_511 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_522 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_533 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_544 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5701__I _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_555 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8082__CLK net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5349__S _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout146_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4385__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4510_ _1180_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout313_I net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5490_ _2133_ mod.Data_Mem.F_M.MRAM\[30\]\[4\] _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4441_ _0642_ mod.Arithmetic.CN.I_in\[51\] _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7363__I mod.Data_Mem.F_M.MRAM\[772\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7160_ _3524_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4372_ _0976_ _1024_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6111_ _1544_ _1506_ _1577_ _2726_ _2727_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _3492_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _2432_ _2658_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6707__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6437__I1 mod.Data_Mem.F_M.MRAM\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout59_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7993_ mod.Instr_Mem.instruction\[30\] net18 net224 mod.Data_Mem.F_M.src\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6944_ _3403_ mod.Data_Mem.F_M.MRAM\[14\]\[6\] _3400_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4073__A1 mod.Arithmetic.CN.I_in\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4073__B2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6875_ mod.Data_Mem.F_M.MRAM\[6\]\[5\] _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8575__CLK net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7538__I _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ mod.Data_Mem.F_M.MRAM\[16\]\[1\] mod.Data_Mem.F_M.MRAM\[17\]\[1\] _2337_ _2450_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5573__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4376__A2 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8545_ _0049_ net327 mod.Data_Mem.F_M.out_data\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5757_ mod.Data_Mem.F_M.MRAM\[770\]\[0\] mod.Data_Mem.F_M.MRAM\[771\]\[0\] _1915_
+ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4708_ _1374_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_159_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8476_ _0572_ net236 mod.Data_Mem.F_M.MRAM\[797\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7314__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5688_ _2277_ _2138_ _2314_ _2316_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_68_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7427_ mod.Data_Mem.F_M.MRAM\[776\]\[6\] _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7273__I mod.Data_Mem.F_M.MRAM\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4639_ _1180_ _1309_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7358_ _3652_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _1978_ _1979_ _1839_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7289_ _3302_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5521__I _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A2 _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4137__I _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4367__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4119__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8448__CLK net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_396 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7559__S _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4047__I mod.Arithmetic.I_out\[72\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6044__A2 mod.Data_Mem.F_M.MRAM\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout263_I net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4990_ _1603_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3941_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6660_ _3220_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5611_ _1747_ mod.Data_Mem.F_M.MRAM\[31\]\[7\] mod.Data_Mem.F_M.MRAM\[30\]\[7\] _2166_
+ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6591_ mod.I_addr\[7\] _3185_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8330_ _0426_ net169 mod.Data_Mem.F_M.MRAM\[777\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5542_ mod.Data_Mem.F_M.MRAM\[797\]\[1\] _2176_ _2177_ mod.Data_Mem.F_M.MRAM\[796\]\[1\]
+ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8261_ _0357_ net92 mod.Data_Mem.F_M.MRAM\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5473_ mod.Data_Mem.F_M.MRAM\[798\]\[1\] mod.Data_Mem.F_M.MRAM\[799\]\[1\] _1880_
+ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7212_ _3564_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5858__A2 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4424_ _0898_ _0984_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8192_ _0302_ net106 mod.Data_Mem.F_M.MRAM\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7143_ _3462_ mod.Data_Mem.F_M.MRAM\[19\]\[7\] _3518_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4355_ _0781_ _0780_ _0800_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__I _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7074_ mod.Data_Mem.F_M.MRAM\[21\]\[0\] _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ _0959_ _0812_ _0875_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6025_ _2641_ mod.Data_Mem.F_M.MRAM\[788\]\[7\] _2642_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5330__I1 mod.Data_Mem.F_M.MRAM\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7607__I0 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ _0202_ net151 mod.Data_Mem.F_M.MRAM\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7965__CLK net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4046__B2 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__C1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6927_ _3392_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout12 net13 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout23 net24 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout34 net36 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6858_ _3351_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout45 net50 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout56 net57 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout67 net68 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5809_ _2209_ mod.Data_Mem.F_M.MRAM\[772\]\[1\] _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5546__A1 mod.Data_Mem.F_M.MRAM\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout78 net96 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4349__A2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout89 net90 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__5546__B2 mod.Data_Mem.F_M.MRAM\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ net6 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8528_ _0032_ net330 mod.Data_Mem.F_M.out_data\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8459_ _0555_ net387 mod.Data_Mem.F_M.MRAM\[795\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5516__I _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6283__S _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5200__B _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6015__C _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8120__CLK net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6810__I mod.Data_Mem.F_M.MRAM\[789\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4760__A2 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5426__I _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4512__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ _0638_ _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout380_I net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6257__I _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _0744_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7988__CLK net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4815__A3 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7830_ _3915_ _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4028__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7761_ _3784_ mod.Data_Mem.F_M.MRAM\[796\]\[7\] _3872_ _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7088__I mod.Data_Mem.F_M.MRAM\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4973_ _1638_ _1640_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6206__B _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6712_ _3258_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7692_ mod.Data_Mem.F_M.MRAM\[792\]\[6\] _3840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6643_ mod.Data_Mem.F_M.MRAM\[25\]\[1\] _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5379__I1 mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6574_ _3173_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4200__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8313_ _0409_ net190 mod.Data_Mem.F_M.MRAM\[775\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5525_ _1815_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4751__A2 mod.Arithmetic.CN.I_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7752__S _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8244_ _0340_ net136 mod.Data_Mem.F_M.MRAM\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5456_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5000__I0 mod.Data_Mem.F_M.MRAM\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4407_ _0721_ _0972_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8175_ mod.DM_en net23 net235 mod.DMen_reg vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5700__A1 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5387_ _2042_ _2048_ _1780_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5700__B2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout202 net204 net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout213 net214 net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7126_ _3433_ _3407_ _3421_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xfanout224 net225 net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout235 net239 net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _0915_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xfanout246 net249 net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_113_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6256__A2 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout257 net258 net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout268 net271 net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_7057_ _3475_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4269_ _0864_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xfanout279 net280 net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6008_ _2400_ mod.Data_Mem.F_M.MRAM\[19\]\[6\] _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7199__S _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6008__A2 mod.Data_Mem.F_M.MRAM\[19\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7056__I1 mod.Data_Mem.F_M.MRAM\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A1 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7959_ _0185_ net322 mod.Data_Mem.F_M.MRAM\[779\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4415__I _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__A2 mod.Arithmetic.CN.I_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__A2 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4258__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6741__S _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout226_I net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6183__A1 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4033__I1 mod.Arithmetic.I_out\[72\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5930__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7572__S _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4060__I mod.Arithmetic.CN.I_in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5310_ _1671_ _1973_ _1884_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6290_ _2053_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5369__S0 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6486__A2 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8164__RN net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _1768_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7371__I mod.Data_Mem.F_M.MRAM\[773\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5172_ _1827_ _1829_ _1834_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_64_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4123_ _0679_ _0682_ _0797_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_96_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4249__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4054_ _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput2 io_in[9] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__8166__CLK net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5997__B2 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__C _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout41_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7813_ mod.Data_Mem.F_M.MRAM\[7\]\[6\] _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7744_ _3230_ _3232_ _3634_ _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _1623_ mod.Data_Mem.F_M.MRAM\[799\]\[0\] _1624_ mod.Data_Mem.F_M.MRAM\[783\]\[0\]
+ _1556_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7675_ _3831_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6626_ _3203_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6174__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6174__B2 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5921__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6557_ _2308_ _2496_ _2662_ _1758_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5508_ _2133_ mod.Data_Mem.F_M.MRAM\[30\]\[7\] _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6488_ _3002_ _3093_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8227_ mod.P1.instr_reg\[9\] net16 net219 mod.P2.dest_reg1\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_79_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8155__RN net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7281__I _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8158_ mod.Data_Mem.F_M.out_data\[68\] net60 net358 mod.Arithmetic.CN.I_in\[68\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6229__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ _3502_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8089_ mod.P2.Rout_reg1\[1\] net35 net261 mod.P2.Rout_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5288__I0 mod.Data_Mem.F_M.MRAM\[773\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5988__A1 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5669__C _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6401__A2 mod.Data_Mem.F_M.MRAM\[781\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A1 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3984__I _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7201__I1 mod.Data_Mem.F_M.MRAM\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__A1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5912__B2 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8146__RN net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6468__A2 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8189__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5140__A2 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5979__B2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout176_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__I0 mod.Data_Mem.F_M.MRAM\[799\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7567__S _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4055__I _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4810_ _1365_ _1382_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_fanout343_I net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _1595_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5600__B1 mod.Data_Mem.F_M.MRAM\[798\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _1208_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6270__I _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7460_ _3703_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4672_ _1338_ _1341_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ _3019_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4706__A2 _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7391_ mod.Data_Mem.F_M.MRAM\[774\]\[4\] _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6342_ _2893_ _2951_ _2952_ _2881_ _1899_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6459__A2 mod.Data_Mem.F_M.MRAM\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8137__RN net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _2842_ _2884_ _2885_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8012_ _0221_ net231 mod.Data_Mem.F_M.MRAM\[14\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5224_ _1609_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5131__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout89_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7259__I1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ _1637_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__A1 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4106_ _0778_ _0779_ _0780_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5086_ mod.Data_Mem.F_M.MRAM\[21\]\[2\] mod.Data_Mem.F_M.MRAM\[20\]\[2\] _1695_ _1753_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4037_ _0688_ mod.Arithmetic.I_out\[74\] _0709_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7187__A3 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5817__S1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5198__A2 _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _2590_ _2009_ _2606_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7727_ _3857_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4939_ _1607_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6147__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7658_ mod.Data_Mem.F_M.MRAM\[790\]\[5\] _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6609_ mod.Data_Mem.F_M.MRAM\[24\]\[0\] _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7589_ _3321_ _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8128__RN net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5524__I _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5122__A2 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A1 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8481__CLK net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3979__I mod.Arithmetic.CN.I_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4076__S _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4633__A1 mod.Arithmetic.CN.I_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6138__A1 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5736__I1 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__B1 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5897__C2 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7489__I1 mod.Data_Mem.F_M.MRAM\[781\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__B2 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout293_I net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7110__I0 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6074__B1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6960_ _3408_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_93_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A1 mod.Arithmetic.CN.I_in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5821__B1 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__C2 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _2378_ _1922_ _2531_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6891_ mod.Data_Mem.F_M.MRAM\[4\]\[5\] _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6377__A1 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5842_ _2157_ mod.Data_Mem.F_M.MRAM\[771\]\[2\] _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8561_ _0065_ net340 mod.Data_Mem.F_M.out_data\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4927__A2 _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6214__B _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5773_ _2396_ _2397_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4513__I _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7512_ _3736_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4724_ _0795_ _1267_ _1269_ _1394_ mod.P3.Res\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8492_ _0588_ net84 mod.Data_Mem.F_M.MRAM\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7443_ mod.Data_Mem.F_M.MRAM\[777\]\[6\] _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4655_ _1223_ _1257_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5727__I1 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7374_ _3660_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4586_ _1220_ _1223_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7629__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6325_ mod.Data_Mem.F_M.MRAM\[13\]\[5\] _2900_ _2901_ mod.Data_Mem.F_M.MRAM\[12\]\[5\]
+ _2936_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6256_ _2868_ _1875_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5104__A2 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5207_ _1555_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6187_ _2177_ _2800_ _2801_ _2710_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5138_ _1580_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5069_ mod.Data_Mem.F_M.MRAM\[6\]\[2\] _1600_ _1644_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6108__C _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7000__S _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4918__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7871__CLK net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6843__A2 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_501 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4854__A1 _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_512 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_523 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_534 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_545 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6056__B1 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_556 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8227__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4082__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4909__A2 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4385__A3 mod.Arithmetic.CN.I_in\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout139_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5365__S _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7644__I mod.Data_Mem.F_M.MRAM\[788\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout306_I net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4440_ mod.Arithmetic.CN.I_in\[52\] _0997_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6531__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5334__A2 _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4371_ _0978_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5164__I _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6110_ _2709_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7090_ mod.Data_Mem.F_M.MRAM\[23\]\[0\] _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7331__I0 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__B1 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _2289_ mod.Data_Mem.F_M.MRAM\[20\]\[7\] _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7992_ mod.Instr_Mem.instruction\[26\] net13 net114 mod.Data_Mem.F_M.src\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6943_ _3255_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4952__B _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6874_ _3359_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ mod.Data_Mem.F_M.MRAM\[14\]\[1\] mod.Data_Mem.F_M.MRAM\[15\]\[1\] _1786_ _2449_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5022__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8544_ _0048_ net327 mod.Data_Mem.F_M.out_data\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5756_ _2099_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5573__A2 mod.Data_Mem.F_M.MRAM\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _1375_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8475_ _0571_ net288 mod.Data_Mem.F_M.MRAM\[797\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5687_ _2315_ mod.Data_Mem.F_M.MRAM\[796\]\[4\] _2280_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7426_ _3686_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6522__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ _0647_ _0958_ _1062_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7894__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7357_ mod.Data_Mem.F_M.MRAM\[772\]\[3\] _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4569_ _1239_ _1131_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ _1976_ _1977_ _1746_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__I0 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7288_ _3608_ _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _2849_ _2852_ _2737_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6834__S _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5249__I _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5693__B _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7561__I0 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6513__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5712__I _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6029__B1 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_397 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout256_I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3940_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6052__I0 mod.Data_Mem.F_M.MRAM\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5610_ _2220_ _2241_ _2244_ _2218_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6590_ _3178_ mod.I_addr\[6\] mod.I_addr\[5\] _3179_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5541_ _2178_ _2180_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8260_ _0356_ net82 mod.Data_Mem.F_M.MRAM\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5472_ _2095_ mod.Data_Mem.F_M.MRAM\[30\]\[1\] _2119_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6211__C _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7211_ _3527_ mod.Data_Mem.F_M.MRAM\[2\]\[1\] _3562_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4423_ _0664_ mod.Arithmetic.CN.I_in\[44\] _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8191_ _0301_ net78 mod.Data_Mem.F_M.MRAM\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7142_ _3521_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4354_ _0942_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7073_ _3483_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4285_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout71_I net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _2526_ mod.Data_Mem.F_M.MRAM\[789\]\[7\] _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8542__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4294__A2 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7607__I1 mod.Data_Mem.F_M.MRAM\[786\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7975_ _0201_ net149 mod.Data_Mem.F_M.MRAM\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6440__B1 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6926_ _3386_ mod.Data_Mem.F_M.MRAM\[14\]\[0\] _3391_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6440__C2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout13 net15 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout24 net39 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6857_ mod.Data_Mem.F_M.MRAM\[779\]\[4\] _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout35 net36 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout57 net66 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5808_ _2389_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout68 net69 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4902__S _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout79 net80 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4349__A3 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _3307_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5546__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8527_ net562 net363 mod.Data_Mem.F_M.out_data\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5739_ _2355_ _2357_ _2358_ _2348_ _2363_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7284__I _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8458_ _0554_ net323 mod.Data_Mem.F_M.MRAM\[795\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6121__C _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7409_ mod.Data_Mem.F_M.MRAM\[775\]\[5\] _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8389_ _0485_ net105 mod.Data_Mem.F_M.MRAM\[785\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5733__S _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8072__CLK net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5857__I0 mod.Data_Mem.F_M.MRAM\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4148__I mod.Arithmetic.CN.I_in\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3987__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6312__B _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7534__I0 _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6739__S _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4767__B _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8565__CLK net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4070_ mod.Arithmetic.I_out\[78\] _0746_ _0709_ mod.Arithmetic.CN.I_in\[22\] _0747_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_77_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout373_I net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7760_ _3875_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ mod.Data_Mem.F_M.MRAM\[5\]\[1\] mod.Data_Mem.F_M.MRAM\[4\]\[1\] _1639_ _1640_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ net10 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7691_ _3839_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5818__S _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6642_ _3211_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5379__I2 mod.Data_Mem.F_M.MRAM\[789\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _3171_ _3172_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4200__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8140__D mod.Data_Mem.F_M.out_data\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8312_ _0408_ net158 mod.Data_Mem.F_M.MRAM\[775\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8095__CLK net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _1844_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4751__A3 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8243_ _0339_ net298 mod.Data_Mem.F_M.MRAM\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5455_ _1496_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4406_ _0620_ _0728_ _0721_ mod.Arithmetic.CN.I_in\[9\] _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_8174_ mod.P2.dest_reg\[8\] net25 net237 mod.Data_Mem.F_M.dest\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5386_ _2008_ _2045_ _2047_ _1833_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5700__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout203 net204 net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout214 net215 net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7125_ _3511_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4337_ _0615_ mod.Arithmetic.ACTI.x\[3\] _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout225 net227 net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout236 net239 net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout247 net248 net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout258 net259 net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7056_ _3462_ mod.Data_Mem.F_M.MRAM\[1\]\[7\] _3465_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout269 net271 net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4268_ _0863_ _0938_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6007_ _2538_ _2624_ _2625_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4199_ mod.Arithmetic.CN.I_in\[24\] _0873_ _0812_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6264__I0 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7958_ _0184_ net382 mod.Data_Mem.F_M.MRAM\[779\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A2 mod.Data_Mem.F_M.MRAM\[789\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6909_ _3246_ mod.Data_Mem.F_M.MRAM\[13\]\[3\] _3376_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7889_ _0115_ net387 mod.Data_Mem.F_M.MRAM\[25\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6911__I _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6192__A2 _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5527__I _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6093__I _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__I0 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout121_I net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4194__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout219_I net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5930__A2 mod.Data_Mem.F_M.MRAM\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5369__S1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5373__S _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5240_ mod.Data_Mem.F_M.MRAM\[773\]\[4\] mod.Data_Mem.F_M.MRAM\[772\]\[4\] _1904_
+ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5694__A1 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6268__I _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _1589_ _1836_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4249__A2 mod.Arithmetic.CN.I_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4053_ mod.Arithmetic.CN.I_in\[12\] _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5997__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6932__S _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7812_ _3904_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7743_ _3865_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout34_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4955_ _1508_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4421__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7674_ mod.Data_Mem.F_M.MRAM\[791\]\[5\] _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4886_ _1553_ _1554_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7746__I0 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6625_ mod.Data_Mem.F_M.MRAM\[26\]\[0\] _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6174__A2 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ _3020_ _2670_ _3157_ _2106_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5507_ _1767_ mod.Data_Mem.F_M.MRAM\[31\]\[7\] _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6487_ _3003_ _2306_ _3026_ _2485_ _2491_ _2499_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_106_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__S _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8226_ _0327_ net242 mod.Data_Mem.F_M.MRAM\[29\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5438_ _1815_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5685__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8157_ mod.Data_Mem.F_M.out_data\[67\] net56 net355 mod.Arithmetic.CN.I_in\[67\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5369_ _2027_ _2028_ _2029_ _2030_ _1896_ _1540_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7108_ _3445_ mod.Data_Mem.F_M.MRAM\[3\]\[0\] _3501_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8088_ mod.P2.Rout_reg1\[0\] net35 net261 mod.P2.Rout_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_48_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5288__I1 mod.Data_Mem.F_M.MRAM\[772\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5437__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7039_ _3464_ _3332_ _3335_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_75_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5810__I _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5988__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7003__S _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8260__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5296__S0 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6165__A2 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4176__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5912__A2 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7472__I _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6088__I _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6752__S _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6779__I1 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5368__S _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4403__A2 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5600__B2 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5595__C _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _1407_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout336_I net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ _1208_ _1210_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6410_ _2369_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7390_ _3668_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ _2011_ _2012_ _1839_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6272_ _1638_ _1907_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8011_ _0220_ net233 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ _1555_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5154_ mod.Data_Mem.F_M.MRAM\[17\]\[3\] mod.Data_Mem.F_M.MRAM\[16\]\[3\] _1543_ _1820_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4105_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4890__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5085_ _1601_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4036_ mod.Arithmetic.CN.I_in\[10\] _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5987_ _2055_ mod.Data_Mem.F_M.MRAM\[786\]\[6\] _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8073__RN net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7726_ mod.Data_Mem.F_M.MRAM\[794\]\[7\] _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4938_ _1574_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _1537_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7657_ _3822_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6147__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7493__S _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6608_ _3194_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7588_ _3783_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6539_ _2571_ mod.Data_Mem.F_M.MRAM\[781\]\[6\] _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7292__I _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8209_ _0310_ net242 mod.Data_Mem.F_M.MRAM\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__S _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4330__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6083__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4633__A2 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5830__A1 _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6386__A2 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4397__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5916__S _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4149__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5897__A1 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5649__A1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4321__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7110__I1 mod.Data_Mem.F_M.MRAM\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6074__A1 mod.Data_Mem.F_M.MRAM\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6074__B2 mod.Data_Mem.F_M.MRAM\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__B1 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5821__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7578__S _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5821__B2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4066__I mod.Arithmetic.CN.I_in\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ _2196_ mod.Data_Mem.F_M.MRAM\[786\]\[4\] _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6890_ _3367_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5841_ _1681_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5098__S _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7377__I mod.Data_Mem.F_M.MRAM\[773\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5772_ mod.Data_Mem.F_M.MRAM\[784\]\[0\] mod.Data_Mem.F_M.MRAM\[785\]\[0\] _1956_
+ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8560_ _0064_ net339 mod.Data_Mem.F_M.out_data\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ _1031_ _1392_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7511_ _3638_ mod.Data_Mem.F_M.MRAM\[782\]\[1\] _3734_ _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8491_ _0587_ net386 mod.Data_Mem.F_M.MRAM\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4015__B mod.Arithmetic.I_out\[72\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5826__S _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7442_ _3694_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4654_ _1286_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7373_ mod.Data_Mem.F_M.MRAM\[773\]\[3\] _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4585_ _1237_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5625__I _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _2902_ _2935_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7629__A2 _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4560__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6688__I0 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6255_ _1581_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6301__A2 _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5206_ _1870_ _1679_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6186_ _1804_ _1734_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5137_ _1731_ _1628_ _1760_ _1762_ _1803_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6456__I _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5068_ _1733_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5812__A1 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4615__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4019_ mod.Arithmetic.I_out\[76\] _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__I _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4379__A1 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _3848_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7317__A1 _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5736__S _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5879__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A2 mod.Data_Mem.F_M.MRAM\[780\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4303__A1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_502 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_513 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_524 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5270__I _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_535 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6056__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_546 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_169_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_557 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__A1 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A1 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__I0 mod.Data_Mem.F_M.MRAM\[771\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5445__I _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6531__A2 mod.Data_Mem.F_M.MRAM\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4370_ _0990_ _1023_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7331__I1 mod.Data_Mem.F_M.MRAM\[771\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A1 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _2320_ mod.Data_Mem.F_M.MRAM\[21\]\[7\] _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6295__B2 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6276__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6047__A1 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__C _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7991_ mod.Instr_Mem.instruction\[24\] net11 net115 mod.Data_Mem.F_M.src\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6942_ _3402_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6873_ mod.Data_Mem.F_M.MRAM\[6\]\[4\] _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5824_ mod.Data_Mem.F_M.MRAM\[30\]\[1\] _1634_ _1921_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5558__B1 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5022__A2 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5755_ _2378_ mod.Data_Mem.F_M.MRAM\[768\]\[0\] _2379_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8543_ _0047_ net251 mod.Data_Mem.F_M.out_data\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ _1242_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5686_ _1649_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8474_ _0570_ net293 mod.Data_Mem.F_M.MRAM\[797\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7425_ mod.Data_Mem.F_M.MRAM\[776\]\[5\] _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4637_ _1178_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8200__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6522__A2 mod.Data_Mem.F_M.MRAM\[768\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7771__S _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7356_ _3651_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4568_ _1126_ _1130_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6307_ _2867_ _2918_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7287_ _3605_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7322__I1 mod.Data_Mem.F_M.MRAM\[770\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4499_ _1055_ _1064_ _1070_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_131_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5333__I0 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6238_ _2850_ _2851_ _2732_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5090__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6169_ _2779_ _2780_ _2781_ _2783_ _2784_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6038__A1 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6119__C _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5958__C _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6210__A1 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7745__I _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6513__A2 mod.Data_Mem.F_M.MRAM\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7561__I1 mod.Data_Mem.F_M.MRAM\[784\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4524__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6277__A1 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5324__I0 mod.Data_Mem.F_M.MRAM\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6029__A1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6029__B2 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8344__CLK net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6824__I mod.Data_Mem.F_M.MRAM\[789\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_398 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6045__B _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4344__I _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout249_I net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8494__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6052__I1 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5376__S _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5540_ _2179_ mod.Data_Mem.F_M.MRAM\[799\]\[1\] mod.Data_Mem.F_M.MRAM\[798\]\[1\]
+ _1917_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4763__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5471_ _1585_ mod.Data_Mem.F_M.MRAM\[31\]\[1\] _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7210_ _3563_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4422_ _1091_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8190_ _0300_ net70 mod.Data_Mem.F_M.MRAM\[19\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7141_ _3460_ mod.Data_Mem.F_M.MRAM\[19\]\[6\] _3518_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4353_ _0945_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_99_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5903__I _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6000__S _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ mod.Data_Mem.F_M.MRAM\[20\]\[7\] _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4284_ mod.Arithmetic.CN.I_in\[27\] _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4818__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _2196_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6935__S _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout64_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7974_ _0200_ net170 mod.Data_Mem.F_M.MRAM\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__A1 _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6440__B2 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6925_ _3390_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_42_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout14 net15 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6856_ _3350_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout25 net38 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout36 net37 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7240__I0 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout47 net49 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout58 net59 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5807_ _2414_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout69 net2 net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3999_ _0654_ _0657_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6787_ mod.Data_Mem.F_M.MRAM\[799\]\[2\] _3306_ _3300_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4754__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8526_ net563 net363 mod.Data_Mem.F_M.out_data\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5738_ _2359_ _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8457_ _0553_ net368 mod.Data_Mem.F_M.MRAM\[795\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5085__I _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5669_ _2296_ mod.Data_Mem.F_M.MRAM\[28\]\[3\] _2298_ _2262_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7408_ _3677_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8388_ _0484_ net104 mod.Data_Mem.F_M.MRAM\[785\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7339_ _3531_ mod.Data_Mem.F_M.MRAM\[771\]\[3\] _3636_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6259__A1 _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__I1 mod.Data_Mem.F_M.MRAM\[17\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6845__S _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6431__A1 _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7231__I0 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7475__I _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4745__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7534__I1 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__A1 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5723__I _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4767__C mod.Arithmetic.ACTI.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7298__I0 _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout199_I net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout366_I net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _1603_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7884__CLK net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ _3257_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7690_ mod.Data_Mem.F_M.MRAM\[792\]\[5\] _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output5_I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6641_ mod.Data_Mem.F_M.MRAM\[25\]\[0\] _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6503__B _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6281__S0 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4736__A1 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _0612_ _3169_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8311_ _0407_ net79 mod.Data_Mem.F_M.MRAM\[774\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5523_ _2131_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6489__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8242_ _0338_ net313 mod.Data_Mem.F_M.MRAM\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5454_ _2076_ _2102_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4405_ _0620_ _0730_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5161__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8173_ mod.P2.dest_reg\[4\] net20 net225 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5385_ _1576_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout204 net213 net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7124_ _3462_ mod.Data_Mem.F_M.MRAM\[3\]\[7\] _3506_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4336_ _0633_ mod.Arithmetic.ACTI.x\[2\] _0846_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout215 net216 net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout226 net227 net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout237 net239 net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7055_ _3474_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout248 net249 net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4267_ _0629_ _0939_ _0941_ mod.P3.Res\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout259 net260 net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_80_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6006_ _2540_ mod.Data_Mem.F_M.MRAM\[21\]\[6\] _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5464__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4198_ mod.Arithmetic.CN.I_in\[26\] _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7957_ _0183_ net231 mod.Data_Mem.F_M.MRAM\[769\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6908_ _3379_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7888_ _0114_ net322 mod.Data_Mem.F_M.MRAM\[25\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7213__I0 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ _3246_ mod.Data_Mem.F_M.MRAM\[769\]\[3\] _3340_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5808__I _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8509_ net572 net357 mod.Data_Mem.F_M.out_data\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5543__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8506__D _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7755__I1 mod.Data_Mem.F_M.MRAM\[796\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4194__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5694__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5170_ mod.Data_Mem.F_M.MRAM\[789\]\[3\] mod.Data_Mem.F_M.MRAM\[788\]\[3\] _1835_
+ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4121_ mod.Arithmetic.ACTI.x\[7\] _0682_ _0795_ mod.Arithmetic.ACTI.x\[6\] _0798_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_111_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4249__A3 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4052_ _0713_ _0714_ _0723_ _0726_ _0727_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_49_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6284__I _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7811_ mod.Data_Mem.F_M.MRAM\[7\]\[5\] _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7742_ mod.Data_Mem.F_M.MRAM\[795\]\[7\] _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8062__CLK net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4954_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout27_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7673_ _3830_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__I _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4885_ _1505_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4709__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6624_ _3202_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5382__A1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _3152_ _3153_ _3154_ _3155_ _3156_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5506_ _2118_ _2146_ _2148_ _2132_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6486_ _2066_ _2497_ _3087_ _3091_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8225_ _0326_ net244 mod.Data_Mem.F_M.MRAM\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5134__A1 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5437_ _2074_ _2071_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5685__A2 mod.Data_Mem.F_M.MRAM\[797\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5368_ mod.Data_Mem.F_M.MRAM\[17\]\[7\] mod.Data_Mem.F_M.MRAM\[16\]\[7\] _1611_ _2030_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8156_ mod.Data_Mem.F_M.out_data\[66\] net58 net357 mod.Arithmetic.CN.I_in\[66\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4893__B1 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ _3500_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4319_ _0929_ _0660_ _0842_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_87_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8087_ _0287_ net81 mod.Data_Mem.F_M.MRAM\[23\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5299_ _1635_ _1961_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5437__A2 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7038_ _3234_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6127__C _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5296__S1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8555__CLK net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5273__I _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A2 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__I mod.Arithmetic.CN.I_in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5600__A2 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout231_I net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4670_ _1339_ _1338_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7922__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout329_I net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5364__A1 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4167__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6561__B1 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5384__S _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6340_ mod.Data_Mem.F_M.MRAM\[789\]\[6\] mod.Data_Mem.F_M.MRAM\[791\]\[6\] mod.Data_Mem.F_M.MRAM\[790\]\[6\]
+ mod.Data_Mem.F_M.MRAM\[788\]\[6\] _2167_ _2315_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6500__C _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6271_ _2868_ _1905_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8010_ _0219_ net305 mod.Data_Mem.F_M.MRAM\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5222_ mod.Data_Mem.F_M.MRAM\[31\]\[4\] _1886_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _1581_ _1818_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4104_ mod.Arithmetic.ACTI.x\[3\] _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ mod.Data_Mem.F_M.MRAM\[22\]\[2\] _1750_ _1644_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4035_ _0681_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8578__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7838__I _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5978__I0 mod.Data_Mem.F_M.MRAM\[784\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _2579_ mod.Data_Mem.F_M.MRAM\[788\]\[6\] _2604_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7592__A2 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7725_ _3856_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4937_ mod.Data_Mem.F_M.MRAM\[790\]\[0\] _1600_ _1602_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7656_ mod.Data_Mem.F_M.MRAM\[790\]\[4\] _3822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4868_ _1527_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ mod.Data_Mem.F_M.MRAM\[11\]\[7\] _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7587_ _3782_ mod.Data_Mem.F_M.MRAM\[785\]\[6\] _3779_ _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4799_ _1315_ _1176_ _1311_ _1468_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _3096_ _2331_ _2623_ _3063_ _3140_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6469_ _2259_ mod.Data_Mem.F_M.MRAM\[13\]\[3\] _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8208_ _0309_ net245 mod.Data_Mem.F_M.MRAM\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8139_ mod.Data_Mem.F_M.out_data\[49\] net53 net331 mod.Arithmetic.CN.I_in\[49\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6083__A2 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5594__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4397__A2 mod.Arithmetic.CN.I_in\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4149__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5897__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4900__I _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5649__A2 mod.Data_Mem.F_M.MRAM\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__I mod.Data_Mem.F_M.dest\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8526__563 net563 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout181_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout279_I net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A3 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A2 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _2457_ _2462_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5771_ _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5178__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7594__S _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7510_ _3735_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4722_ _1270_ _1391_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8490_ _0586_ net145 mod.Data_Mem.F_M.MRAM\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7441_ mod.Data_Mem.F_M.MRAM\[777\]\[5\] _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8100__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4653_ _1287_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7372_ _3659_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4584_ _1238_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6323_ _2903_ mod.Data_Mem.F_M.MRAM\[15\]\[5\] mod.Data_Mem.F_M.MRAM\[14\]\[5\] _2253_
+ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4560__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6688__I1 mod.Data_Mem.F_M.MRAM\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _2679_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout94_I net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ mod.Data_Mem.F_M.MRAM\[15\]\[4\] _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__I _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6185_ _2325_ mod.Data_Mem.F_M.MRAM\[6\]\[2\] mod.Data_Mem.F_M.MRAM\[7\]\[2\] _2753_
+ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _1782_ _1802_ _1676_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7769__S _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ mod.Data_Mem.F_M.MRAM\[5\]\[2\] mod.Data_Mem.F_M.MRAM\[4\]\[2\] _1639_ _1734_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4018_ _0686_ _0687_ _0688_ _0689_ _0692_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_4
XANTENNA__5289__S _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6405__C _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4379__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ _2391_ mod.Data_Mem.F_M.MRAM\[782\]\[5\] _2588_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7708_ mod.Data_Mem.F_M.MRAM\[793\]\[6\] _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4921__S _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7317__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5328__A1 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7639_ _3813_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7009__S _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5816__I _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5879__A2 mod.Data_Mem.F_M.MRAM\[771\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5752__S _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4303__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5500__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_503 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_514 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_525 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_536 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_547 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_558 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5500__B _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8514__D _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7556__A2 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4790__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5726__I _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4542__A2 mod.Arithmetic.CN.I_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A2 mod.Data_Mem.F_M.MRAM\[783\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4077__I mod.Arithmetic.ACTI.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6047__A2 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7990_ mod.Instr_Mem.instruction\[23\] net11 net100 mod.Data_Mem.F_M.src\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ _3253_ mod.Data_Mem.F_M.MRAM\[14\]\[5\] _3400_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6872_ _3358_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5558__A1 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5823_ _2359_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5558__B2 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8542_ _0046_ net253 mod.Data_Mem.F_M.out_data\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5754_ _1717_ mod.Data_Mem.F_M.MRAM\[769\]\[0\] _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ _0646_ mod.Arithmetic.ACTI.x\[6\] _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4781__A2 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8473_ _0569_ net291 mod.Data_Mem.F_M.MRAM\[797\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5636__I _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5685_ _2128_ mod.Data_Mem.F_M.MRAM\[797\]\[4\] _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7424_ _3685_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4636_ _1058_ _1305_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7355_ mod.Data_Mem.F_M.MRAM\[772\]\[2\] _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4567_ _0664_ mod.Arithmetic.CN.I_in\[68\] _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_78_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6306_ _2914_ _2915_ _2916_ _2917_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7286_ _3607_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _1069_ _1071_ _1068_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6237_ _1577_ _1857_ _2727_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4297__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5494__B1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6168_ _2678_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7499__S _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5119_ _1649_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ _2713_ _2714_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8146__CLK net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5341__S0 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__A1 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6135__C _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5549__A1 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8296__CLK net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__I0 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4524__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6277__A2 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5324__I1 mod.Data_Mem.F_M.MRAM\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6029__A2 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5788__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_399 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4460__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6201__A2 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout144_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5960__A1 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5456__I _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout311_I net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _2086_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8194__RN net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4421_ _1092_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8019__CLK net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7140_ _3520_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4352_ _0948_ _1025_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6287__I _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7071_ _3482_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5315__I1 mod.Data_Mem.F_M.MRAM\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4283_ _0877_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4279__A1 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4818__A3 mod.Arithmetic.I_out\[79\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6022_ _2622_ _2640_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8169__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7112__S _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7973_ _0199_ net72 mod.Data_Mem.F_M.MRAM\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout57_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__I _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6924_ _3235_ _3387_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6440__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6855_ mod.Data_Mem.F_M.MRAM\[779\]\[3\] _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout15 net24 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout26 net33 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout37 net38 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7240__I1 mod.Data_Mem.F_M.MRAM\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5806_ mod.Data_Mem.F_M.MRAM\[782\]\[1\] mod.Data_Mem.F_M.MRAM\[783\]\[1\] _1711_
+ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout59 net65 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4203__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6786_ _3305_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3998_ _0660_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8525_ net564 net357 mod.Data_Mem.F_M.out_data\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5737_ _2360_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4754__A2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8456_ _0552_ net317 mod.Data_Mem.F_M.MRAM\[795\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _2297_ _2206_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7407_ mod.Data_Mem.F_M.MRAM\[775\]\[4\] _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5703__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4619_ _1288_ _0730_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7581__I _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8387_ _0483_ net180 mod.Data_Mem.F_M.MRAM\[785\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5599_ mod.Data_Mem.F_M.MRAM\[29\]\[5\] _2221_ _2222_ mod.Data_Mem.F_M.MRAM\[28\]\[5\]
+ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_85_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7338_ _3641_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6259__A2 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7269_ mod.Data_Mem.F_M.MRAM\[5\]\[2\] _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6925__I _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A2 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5477__S _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7231__I1 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6195__A1 _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5942__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4745__A2 mod.Arithmetic.CN.I_in\[71\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8176__RN net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6498__A2 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7298__I1 mod.Data_Mem.F_M.MRAM\[768\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4681__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8461__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout261_I net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7470__I1 mod.Data_Mem.F_M.MRAM\[780\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout359_I net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4970_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _3210_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6186__A1 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6571_ mod.I_addr\[2\] _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5933__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6281__S1 _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8310_ _0406_ net85 mod.Data_Mem.F_M.MRAM\[774\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5522_ _2076_ _2061_ _2155_ _2161_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8241_ _0337_ net312 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5453_ _2098_ _2101_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5914__I _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4404_ _1049_ _1075_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8172_ mod.P2.dest_reg\[2\] net21 net225 mod.Data_Mem.F_M.dest\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_132_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5384_ mod.Data_Mem.F_M.MRAM\[785\]\[7\] mod.Data_Mem.F_M.MRAM\[784\]\[7\] _1889_
+ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5161__A2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7123_ _3510_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout205 net208 net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4335_ mod.Arithmetic.CN.I_in\[64\] _0918_ mod.Arithmetic.ACTI.x\[1\] _0634_ _1009_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_59_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout216 net217 net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout227 net228 net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout238 net239 net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7054_ _3460_ mod.Data_Mem.F_M.MRAM\[1\]\[6\] _3469_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout249 net250 net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4266_ _0774_ _0857_ _0859_ _0940_ _0627_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4121__B1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6745__I _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6005_ _2259_ mod.Data_Mem.F_M.MRAM\[20\]\[6\] _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4197_ _0637_ _0811_ _0871_ _0814_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7956_ _0182_ net135 mod.Data_Mem.F_M.MRAM\[769\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6907_ _3243_ mod.Data_Mem.F_M.MRAM\[13\]\[2\] _3376_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7887_ _0113_ net157 mod.Data_Mem.F_M.MRAM\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7213__I1 mod.Data_Mem.F_M.MRAM\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6838_ _3341_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6177__A1 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5924__A1 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _3291_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5096__I _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8508_ net573 net359 mod.Data_Mem.F_M.out_data\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8439_ _0535_ net373 mod.Data_Mem.F_M.MRAM\[792\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8484__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6101__A1 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4663__A1 mod.Arithmetic.CN.I_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7486__I _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5000__S _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4718__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout107_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5694__A3 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4120_ _0789_ _0793_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_122_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4051_ mod.Arithmetic.CN.I_in\[11\] _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_96_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7810_ _3903_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _3864_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4953_ _1500_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6514__B _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7672_ mod.Data_Mem.F_M.MRAM\[791\]\[4\] _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4884_ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6623_ mod.Data_Mem.F_M.MRAM\[24\]\[7\] _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5906__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6954__I0 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5757__I1 mod.Data_Mem.F_M.MRAM\[771\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6554_ _2538_ _2666_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5382__A2 mod.Data_Mem.F_M.MRAM\[786\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5505_ _1783_ mod.Data_Mem.F_M.MRAM\[798\]\[6\] _2147_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6485_ _3026_ _2502_ _3090_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8224_ _0325_ net248 mod.Data_Mem.F_M.MRAM\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _2066_ _2068_ _2070_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5134__A2 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8155_ mod.Data_Mem.F_M.out_data\[65\] net56 net336 mod.Arithmetic.CN.I_in\[65\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5367_ mod.Data_Mem.F_M.MRAM\[19\]\[7\] mod.Data_Mem.F_M.MRAM\[18\]\[7\] _1809_ _2029_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4893__A1 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7106_ _3433_ _3272_ _3407_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4893__B2 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4318_ _0911_ _0991_ _0927_ _0933_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8086_ _0286_ net78 mod.Data_Mem.F_M.MRAM\[23\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5298_ mod.Data_Mem.F_M.MRAM\[783\]\[5\] _1934_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7037_ _3463_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4249_ _0655_ mod.Arithmetic.CN.I_in\[57\] _0663_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__A1 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3999__A3 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6398__A1 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7300__S _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7939_ _0165_ net100 mod.Data_Mem.F_M.MRAM\[799\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4176__A3 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4581__B1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5554__I _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7122__I0 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__I0 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout224_I net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__A1 mod.Data_Mem.F_M.MRAM\[781\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6561__B2 mod.Data_Mem.F_M.MRAM\[769\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6270_ _2679_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _1678_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5152_ mod.Data_Mem.F_M.MRAM\[19\]\[3\] mod.Data_Mem.F_M.MRAM\[18\]\[3\] _1651_ _1818_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6077__B1 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4103_ mod.Arithmetic.CN.I_in\[11\] _0727_ _0752_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5083_ _1599_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4627__A1 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4034_ _0680_ mod.Arithmetic.I_out\[79\] _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7120__S _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5978__I1 mod.Data_Mem.F_M.MRAM\[785\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5985_ _2464_ mod.Data_Mem.F_M.MRAM\[789\]\[6\] _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6244__B _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5052__A1 _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5639__I _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7724_ mod.Data_Mem.F_M.MRAM\[794\]\[6\] _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4936_ mod.Data_Mem.F_M.MRAM\[789\]\[0\] mod.Data_Mem.F_M.MRAM\[788\]\[0\] _1604_
+ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7655_ _3821_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4867_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6606_ _3193_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7586_ _3318_ _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6552__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4798_ _1315_ _1176_ _1311_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6537_ _2065_ _2496_ _2628_ _1758_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_119_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7790__S _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6304__A1 _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6468_ _3016_ mod.Data_Mem.F_M.MRAM\[1\]\[3\] _2635_ _3073_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8207_ _0308_ net243 mod.Data_Mem.F_M.MRAM\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ _2075_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6399_ _2487_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8138_ mod.Data_Mem.F_M.out_data\[48\] net59 net348 mod.Arithmetic.CN.I_in\[48\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8069_ _0278_ net75 mod.Data_Mem.F_M.MRAM\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7030__S _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8072__D mod.P3.Res\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6918__I0 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7764__I _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6543__A1 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7205__S _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8052__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4321__A3 mod.Arithmetic.CN.I_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6059__B1 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5233__B _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4085__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5282__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6064__B _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout341_I net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5770_ _2087_ _1553_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4721_ _1270_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6909__I0 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7440_ _3693_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ _1298_ _1301_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7582__I0 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7371_ mod.Data_Mem.F_M.MRAM\[773\]\[2\] _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4583_ _1250_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6322_ _2919_ _2922_ _2929_ _2933_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7334__I0 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _2865_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__I0 mod.Data_Mem.F_M.MRAM\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5204_ _1805_ _1806_ _1869_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout87_I net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6184_ _2794_ _2798_ _2696_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6239__B _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6954__S _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5135_ _1598_ _1800_ _1801_ _1561_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _1732_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4017_ _0693_ mod.Arithmetic.I_out\[74\] _0690_ mod.Arithmetic.I_out\[73\] _0694_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_38_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5968_ _1774_ mod.Data_Mem.F_M.MRAM\[783\]\[5\] _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7707_ _3847_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4919_ _1567_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5981__C1 _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5899_ _2447_ _2519_ _2520_ _2219_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5328__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6525__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7638_ mod.Data_Mem.F_M.MRAM\[788\]\[3\] _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7569_ _3292_ _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8075__CLK net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6928__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5500__A2 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_504 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_515 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_526 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7912__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_537 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_548 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_559 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__B1 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5016__A1 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7308__A3 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8530__D _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5742__I _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout291_I net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout389_I net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _3401_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6871_ mod.Data_Mem.F_M.MRAM\[6\]\[3\] _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5822_ _2346_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5558__A2 mod.Data_Mem.F_M.MRAM\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5753_ _2142_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8541_ _0045_ net271 mod.Data_Mem.F_M.out_data\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5917__I _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8098__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4821__I _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _0641_ mod.Arithmetic.ACTI.x\[5\] _1125_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6507__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8472_ _0568_ net287 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5684_ _2308_ _2135_ _2310_ _2312_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7423_ mod.Data_Mem.F_M.MRAM\[776\]\[4\] _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4635_ _1170_ _1171_ _1180_ _1181_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_159_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5853__S _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7354_ _3650_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _1124_ _1132_ _1133_ _1138_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6305_ _2873_ _1970_ _2782_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7285_ _3603_ mod.Data_Mem.F_M.MRAM\[768\]\[0\] _3606_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4497_ _1053_ _1167_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6236_ _2156_ _1853_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4297__A2 mod.Arithmetic.CN.I_in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5494__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5494__B2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6684__S _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6167_ _1737_ _1688_ _2782_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5118_ _1783_ mod.Data_Mem.F_M.MRAM\[791\]\[2\] _1784_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6098_ _1830_ _1590_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5049_ _1704_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5341__S1 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5797__A2 mod.Data_Mem.F_M.MRAM\[789\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7546__I0 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3980__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4524__A3 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A1 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6393__I _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4906__I _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__A2 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4460__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5960__A2 mod.Data_Mem.F_M.MRAM\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout304_I net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4420_ _0834_ mod.Arithmetic.CN.I_in\[35\] _0830_ _0893_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4515__A3 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4351_ _0951_ _0976_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7070_ mod.Data_Mem.F_M.MRAM\[20\]\[6\] _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4282_ _0667_ mod.Arithmetic.CN.I_in\[19\] _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4279__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6021_ _1676_ _2117_ _2631_ _2639_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_98_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7972_ _0198_ net80 mod.Data_Mem.F_M.MRAM\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6923_ _3388_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6854_ _3349_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7776__I0 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout16 net18 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout27 net33 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout38 net39 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_50_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5805_ _2427_ _1713_ _2428_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6785_ net5 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4203__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3997_ _0663_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8524_ net565 net357 mod.Data_Mem.F_M.out_data\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5736_ mod.Data_Mem.F_M.MRAM\[2\]\[0\] mod.Data_Mem.F_M.MRAM\[3\]\[0\] _1971_ _2361_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7528__I0 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8455_ _0551_ net369 mod.Data_Mem.F_M.MRAM\[794\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5667_ _1611_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ mod.Arithmetic.CN.I_in\[14\] _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7406_ _3676_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8386_ _0482_ net181 mod.Data_Mem.F_M.MRAM\[785\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ _2223_ _2233_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5703__A2 mod.Data_Mem.F_M.MRAM\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7337_ _3640_ mod.Data_Mem.F_M.MRAM\[771\]\[2\] _3636_ _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6478__I _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4549_ _1122_ _1139_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7268_ _3596_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8113__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6219_ _2709_ _2678_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7199_ _3533_ mod.Data_Mem.F_M.MRAM\[29\]\[4\] _3553_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7303__S _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8263__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A2 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__S _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7767__I0 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A2 mod.Data_Mem.F_M.MRAM\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4461__I mod.Arithmetic.CN.I_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7772__I _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5292__I _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5458__A1 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7213__S _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4681__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5630__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout254_I net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5467__I _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4197__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6570_ _3170_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5933__A2 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5521_ _2112_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8240_ _0336_ net298 mod.Data_Mem.F_M.MRAM\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5452_ _2100_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4403_ _0894_ _0832_ _0980_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_126_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8171_ mod.P2.dest_reg\[1\] net21 net227 mod.Data_Mem.F_M.dest\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5383_ _1767_ _2043_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7122_ _3460_ mod.Data_Mem.F_M.MRAM\[3\]\[6\] _3506_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4334_ _0646_ mod.Arithmetic.CN.I_in\[67\] _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5135__C _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout206 net208 net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout217 net393 net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout228 net234 net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7053_ _1968_ _3466_ _3473_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout239 net240 net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4265_ _0774_ _0779_ _0800_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4121__A1 mod.Arithmetic.ACTI.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6004_ mod.Data_Mem.F_M.MRAM\[16\]\[6\] mod.Data_Mem.F_M.MRAM\[17\]\[6\] _1937_ _2623_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4121__B2 mod.Arithmetic.ACTI.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4196_ _0645_ _0810_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7955_ _0181_ net122 mod.Data_Mem.F_M.MRAM\[769\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6906_ _3378_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7886_ _0112_ net386 mod.Data_Mem.F_M.MRAM\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _3243_ mod.Data_Mem.F_M.MRAM\[769\]\[2\] _3340_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7793__S _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6768_ mod.Data_Mem.F_M.MRAM\[8\]\[7\] _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8507_ _0011_ net345 mod.Data_Mem.F_M.out_data\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5719_ _2344_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6699_ _3248_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8438_ _0534_ net379 mod.Data_Mem.F_M.MRAM\[792\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5688__A1 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5232__S0 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8369_ _0465_ net291 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6101__A2 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7033__S _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4112__B2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5061__B _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8075__D mod.P3.Res\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8094__RN net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5612__A1 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8009__CLK net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__I0 mod.Data_Mem.F_M.MRAM\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5750__I _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__I0 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ _0686_ mod.Arithmetic.I_out\[75\] _0719_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5603__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5603__B2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7740_ mod.Data_Mem.F_M.MRAM\[795\]\[6\] _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4952_ _1579_ _1593_ _1598_ _1620_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_17_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5197__I _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7671_ _3829_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4883_ mod.Data_Mem.F_M.src\[2\] _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6159__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6622_ _3201_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5906__A2 mod.Data_Mem.F_M.MRAM\[789\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6954__I1 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6553_ _2722_ mod.Data_Mem.F_M.MRAM\[13\]\[7\] _2387_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5504_ _1615_ mod.Data_Mem.F_M.MRAM\[799\]\[6\] _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6484_ _2431_ _3088_ _3089_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8223_ _0324_ net244 mod.Data_Mem.F_M.MRAM\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5435_ _2086_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6331__A2 _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4342__A1 _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ mod.Data_Mem.F_M.MRAM\[21\]\[7\] mod.Data_Mem.F_M.MRAM\[20\]\[7\] _1880_ _2028_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8154_ mod.Data_Mem.F_M.out_data\[64\] net60 net348 mod.Arithmetic.CN.I_in\[64\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4893__A2 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7105_ _3499_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4317_ _0921_ _0926_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8085_ _0285_ net88 mod.Data_Mem.F_M.MRAM\[23\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5297_ _1888_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7036_ _3462_ mod.Data_Mem.F_M.MRAM\[18\]\[7\] _3457_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7831__A2 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4248_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7788__S _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4645__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5842__A1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6692__S _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4179_ _0807_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_67_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8076__RN net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6491__I _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7938_ _0164_ net97 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7869_ _0095_ net320 mod.Data_Mem.F_M.MRAM\[11\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7028__S _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4581__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4581__B2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4333__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7122__I1 mod.Data_Mem.F_M.MRAM\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6086__A1 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5133__I0 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5833__A1 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8533__D _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4914__I _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5597__B1 mod.Data_Mem.F_M.MRAM\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__I1 mod.Data_Mem.F_M.MRAM\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__C1 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4021__B1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6561__A2 _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4572__A1 mod.Arithmetic.CN.I_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout217_I net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5220_ _1872_ _1883_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4324__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4324__B2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ mod.Data_Mem.F_M.MRAM\[3\]\[3\] mod.Data_Mem.F_M.MRAM\[1\]\[3\] mod.Data_Mem.F_M.MRAM\[0\]\[3\]
+ mod.Data_Mem.F_M.MRAM\[2\]\[3\] _1816_ _1787_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6077__A1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4102_ _0760_ _0772_ _0773_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6077__B2 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5082_ _1746_ _1748_ _1565_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4033_ _0637_ mod.Arithmetic.I_out\[72\] _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8324__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__S _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _2550_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5052__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6244__C _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout32_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7723_ _3855_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4935_ _1603_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_75_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5856__S _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7654_ mod.Data_Mem.F_M.MRAM\[790\]\[3\] _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4866_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6001__A1 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6605_ mod.Data_Mem.F_M.MRAM\[11\]\[6\] _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7585_ _3781_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6552__A2 mod.Data_Mem.F_M.MRAM\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ _1313_ _1317_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6536_ _3013_ _3134_ _3138_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6304__A2 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6467_ _2169_ mod.Data_Mem.F_M.MRAM\[0\]\[3\] _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8206_ _0307_ net299 mod.Data_Mem.F_M.MRAM\[12\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5418_ _1511_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6398_ _3002_ _3006_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5349_ mod.Data_Mem.F_M.MRAM\[785\]\[6\] mod.Data_Mem.F_M.MRAM\[784\]\[6\] _1889_
+ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8137_ mod.Data_Mem.F_M.out_data\[47\] net44 net255 mod.Arithmetic.CN.I_in\[47\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8068_ _0277_ net91 mod.Data_Mem.F_M.MRAM\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5815__A1 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ _3451_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5579__B1 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6918__I1 mod.Data_Mem.F_M.MRAM\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4306__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8528__D _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6059__A1 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6059__B2 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__S _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5282__A2 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7020__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8497__CLK net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6231__A1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _1273_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4793__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout334_I net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5990__B1 _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__I1 mod.Data_Mem.F_M.MRAM\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _1303_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6080__B _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7582__I1 mod.Data_Mem.F_M.MRAM\[785\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4545__A1 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7370_ _3658_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ _1018_ _1251_ _1136_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6321_ _2879_ _2931_ _2932_ _2897_ _1675_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7334__I1 mod.Data_Mem.F_M.MRAM\[771\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6252_ _2695_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5203_ _1632_ _1862_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5896__I1 mod.Data_Mem.F_M.MRAM\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6183_ _2680_ _2797_ _2693_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5134_ mod.Data_Mem.F_M.MRAM\[799\]\[2\] _1780_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6845__I0 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5065_ _1567_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6470__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4016_ _0688_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_38_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4554__I mod.Arithmetic.CN.I_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5967_ _2520_ _2578_ _2586_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6773__A2 mod.Data_Mem.F_M.dest\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7706_ mod.Data_Mem.F_M.MRAM\[793\]\[5\] _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4784__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4918_ _1582_ _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5981__B1 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5898_ _2116_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7637_ _3812_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6525__A2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4849_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7568_ _3770_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6519_ _3120_ _3122_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7499_ _3645_ mod.Data_Mem.F_M.MRAM\[781\]\[5\] _3726_ _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7306__S _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5334__B _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_505 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_516 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_527 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_538 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__S _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_549 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6461__A1 mod.Data_Mem.F_M.MRAM\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4862__I2 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5016__A2 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7261__I0 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__A1 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout284_I net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7887__CLK net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6870_ _3357_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6204__A1 _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7252__I0 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5821_ _2440_ _2441_ _2442_ _2360_ _2443_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_62_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8540_ _0044_ net269 mod.Data_Mem.F_M.out_data\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4766__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ mod.Data_Mem.F_M.MRAM\[782\]\[0\] mod.Data_Mem.F_M.MRAM\[783\]\[0\] _2376_
+ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4703_ mod.Arithmetic.CN.I_in\[67\] _1246_ _0642_ mod.Arithmetic.ACTI.x\[4\] _1374_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8471_ _0567_ net238 mod.Data_Mem.F_M.MRAM\[796\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5683_ _2169_ mod.Data_Mem.F_M.MRAM\[28\]\[4\] _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7422_ _3684_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4634_ _1180_ _1181_ _1170_ _1171_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7353_ mod.Data_Mem.F_M.MRAM\[772\]\[1\] _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5191__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4565_ _1235_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6304_ _2855_ _1972_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7284_ _3605_ _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4496_ _1054_ _1056_ _1067_ _1072_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6235_ _2842_ _2847_ _2848_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__I3 _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5494__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ _2708_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _1658_ mod.Data_Mem.F_M.MRAM\[790\]\[2\] _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6097_ _2008_ _1586_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ _1648_ _1715_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4284__I mod.Arithmetic.CN.I_in\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _3438_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4757__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7546__I1 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3980__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__S _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6131__B1 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__A2 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6674__I _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__A1 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7482__I0 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8541__D _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4922__I _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4748__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6342__C _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5753__I _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4350_ _0978_ _0990_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4281_ _0879_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6020_ _2372_ _2634_ _2638_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7473__I0 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7971_ _0197_ net158 mod.Data_Mem.F_M.MRAM\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6922_ mod.Data_Mem.F_M.dest\[1\] _3333_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__I0 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ mod.Data_Mem.F_M.MRAM\[779\]\[2\] _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7776__I1 mod.Data_Mem.F_M.MRAM\[797\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout17 net18 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4832__I mod.Data_Mem.F_M.src\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout28 net29 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4739__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5804_ _1791_ mod.Data_Mem.F_M.MRAM\[771\]\[1\] _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout39 net69 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6784_ _3304_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3996_ _0666_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8523_ _0027_ net355 mod.Data_Mem.F_M.out_data\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5735_ _2349_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7528__I1 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8454_ _0550_ net168 mod.Data_Mem.F_M.MRAM\[794\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7902__CLK net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5666_ _1787_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7405_ mod.Data_Mem.F_M.MRAM\[775\]\[3\] _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4617_ mod.Arithmetic.CN.I_in\[13\] _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8385_ _0481_ net181 mod.Data_Mem.F_M.MRAM\[785\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5597_ _2224_ mod.Data_Mem.F_M.MRAM\[31\]\[5\] mod.Data_Mem.F_M.MRAM\[30\]\[5\] _2225_
+ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_85_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7336_ _3305_ _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _1205_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7267_ mod.Data_Mem.F_M.MRAM\[5\]\[1\] _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4479_ _1044_ _1045_ _1143_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6218_ _1614_ _1820_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7198_ _2206_ _3550_ _3556_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ _2582_ mod.Data_Mem.F_M.MRAM\[22\]\[1\] mod.Data_Mem.F_M.MRAM\[23\]\[1\] _2753_
+ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6416__A1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4943__S _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8558__CLK net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7767__I1 mod.Data_Mem.F_M.MRAM\[797\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6162__C _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5155__A1 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8088__CLK net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__S _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A2 mod.Data_Mem.F_M.MRAM\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7925__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ mod.Data_Mem.F_M.MRAM\[29\]\[0\] _2083_ _2156_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5451_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4402_ _1052_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8170_ mod.P2.dest_reg\[0\] net20 net223 mod.Data_Mem.F_M.dest\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5382_ _1923_ mod.Data_Mem.F_M.MRAM\[786\]\[7\] _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7121_ _3509_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4333_ _0915_ _1005_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout207 net212 net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout218 net220 net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout229 net231 net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_7052_ _3316_ _3466_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4264_ _0863_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_86_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5854__C1 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _2409_ _2610_ _2616_ _2618_ _2621_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_132_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4827__I mod.Data_Mem.F_M.src\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4195_ _0638_ _0815_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7954_ _0180_ net135 mod.Data_Mem.F_M.MRAM\[769\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6905_ _3240_ mod.Data_Mem.F_M.MRAM\[13\]\[1\] _3376_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7885_ _0111_ net379 mod.Data_Mem.F_M.MRAM\[26\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6836_ _3336_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_62_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5385__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _3290_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3979_ mod.Arithmetic.CN.I_in\[40\] _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ _0010_ net348 mod.Data_Mem.F_M.out_data\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5718_ _2062_ _2340_ _2343_ _2164_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6698_ net7 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7126__A2 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5137__A1 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8437_ _0533_ net192 mod.Data_Mem.F_M.MRAM\[792\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5393__I _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5137__B2 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5649_ _2157_ mod.Data_Mem.F_M.MRAM\[28\]\[1\] _2280_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5688__A2 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5232__S1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8368_ _0464_ net287 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7319_ _1851_ _3626_ _3629_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8299_ _0395_ net143 mod.Data_Mem.F_M.MRAM\[773\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__B _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8380__CLK net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6412__I1 mod.Data_Mem.F_M.MRAM\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7783__I _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6399__I _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5128__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5236__C _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5300__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7023__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout197_I net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5151__I1 mod.Data_Mem.F_M.MRAM\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7053__A1 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A3 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _1566_ _1606_ _1613_ _1618_ _1619_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_36_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output3_I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7670_ mod.Data_Mem.F_M.MRAM\[791\]\[3\] _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4882_ _1509_ _1531_ _1532_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6621_ mod.Data_Mem.F_M.MRAM\[24\]\[6\] _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8103__CLK net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__B1 _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6552_ _2410_ mod.Data_Mem.F_M.MRAM\[12\]\[7\] _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5503_ _2133_ mod.Data_Mem.F_M.MRAM\[30\]\[6\] _2145_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_9_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6483_ _2526_ mod.Data_Mem.F_M.MRAM\[780\]\[3\] _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8222_ _0323_ net311 mod.Data_Mem.F_M.MRAM\[29\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5434_ _2085_ _2061_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A2 _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8153_ mod.Data_Mem.F_M.out_data\[63\] net61 net361 mod.Arithmetic.CN.I_in\[63\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5365_ mod.Data_Mem.F_M.MRAM\[23\]\[7\] mod.Data_Mem.F_M.MRAM\[22\]\[7\] _1878_ _2027_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5941__I _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7104_ mod.Data_Mem.F_M.MRAM\[23\]\[7\] _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4316_ _0988_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8084_ _0284_ net73 mod.Data_Mem.F_M.MRAM\[23\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6258__B _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5296_ _1952_ _1953_ _1958_ _1959_ _1882_ _1645_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5827__C1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6095__A2 _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ _3258_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4247_ mod.Arithmetic.CN.I_in\[58\] _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__A2 mod.Data_Mem.F_M.MRAM\[771\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _0823_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7937_ _0163_ net288 mod.Data_Mem.F_M.MRAM\[799\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7868_ _0094_ net378 mod.Data_Mem.F_M.MRAM\[11\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6819_ _3328_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7799_ _3322_ mod.Data_Mem.F_M.MRAM\[798\]\[7\] _3894_ _3898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4030__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5530__A1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7283__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6086__A2 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__I1 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5833__A2 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5597__A1 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8126__CLK net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__B2 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6546__B1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6546__C2 _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__A2 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4930__I _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4572__A2 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout112_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4324__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5150_ _1815_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4101_ _0774_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6077__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ mod.Data_Mem.F_M.MRAM\[19\]\[2\] mod.Data_Mem.F_M.MRAM\[18\]\[2\] _1747_ _1748_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4032_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5983_ _2407_ _2587_ _2602_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7722_ mod.Data_Mem.F_M.MRAM\[794\]\[5\] _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4934_ _1517_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7329__A2 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7653_ _3820_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout25_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4865_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5936__I _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6001__A2 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4840__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6604_ _3192_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _3754_ mod.Data_Mem.F_M.MRAM\[785\]\[5\] _3779_ _3781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4796_ _1303_ _1321_ _1465_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6968__S _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6535_ _3059_ _2636_ _2637_ _3019_ _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5760__A1 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6466_ _3062_ _3072_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8205_ _0306_ net297 mod.Data_Mem.F_M.MRAM\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5417_ _2074_ _2071_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6397_ _3003_ _2256_ _3004_ _2401_ _2397_ _3005_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8136_ mod.Data_Mem.F_M.out_data\[46\] net44 net251 mod.Arithmetic.CN.I_in\[46\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5348_ _1921_ _2009_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7799__S _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8067_ _0276_ net82 mod.Data_Mem.F_M.MRAM\[21\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5279_ _1936_ _1940_ _1942_ _1566_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7018_ _3450_ mod.Data_Mem.F_M.MRAM\[18\]\[1\] _3448_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A1 mod.Data_Mem.F_M.MRAM\[797\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6379__I0 mod.Data_Mem.F_M.MRAM\[789\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4306__A2 mod.Arithmetic.CN.I_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__A2 mod.Data_Mem.F_M.MRAM\[782\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7502__S _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__S0 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout390 net391 net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__8544__D _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6231__A2 _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5990__A1 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4793__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5756__I _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5990__B2 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4660__I mod.Arithmetic.CN.I_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4650_ _1304_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_fanout327_I net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _1252_ _1251_ _1136_ _1017_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6320_ _1945_ _1947_ _2895_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6251_ _2367_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5202_ _1864_ _1866_ _1867_ _1702_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6182_ mod.Data_Mem.F_M.MRAM\[13\]\[2\] _2193_ _1813_ mod.Data_Mem.F_M.MRAM\[12\]\[2\]
+ _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_111_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5133_ _1785_ _1790_ _1795_ _1799_ _1526_ _1530_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5064_ _1538_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4015_ _0690_ mod.Arithmetic.I_out\[73\] mod.Arithmetic.I_out\[72\] _0691_ _0692_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__4835__I mod.Data_Mem.F_M.src\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8441__CLK net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5867__S _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _2557_ _2581_ _2585_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5281__I0 mod.Data_Mem.F_M.MRAM\[787\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7705_ _3846_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4917_ mod.Data_Mem.F_M.MRAM\[771\]\[0\] mod.Data_Mem.F_M.MRAM\[770\]\[0\] _1585_
+ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5981__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8591__CLK net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5666__I _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _2126_ _2348_ _2350_ _2517_ _2518_ _2355_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5981__B2 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7636_ mod.Data_Mem.F_M.MRAM\[788\]\[2\] _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _1503_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7567_ _3731_ mod.Data_Mem.F_M.MRAM\[784\]\[7\] _3759_ _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4779_ _1307_ _1319_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6518_ _2827_ _3121_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7498_ _3727_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6449_ _2320_ mod.Data_Mem.F_M.MRAM\[769\]\[2\] _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8119_ mod.Data_Mem.F_M.out_data\[29\] net43 net278 mod.Arithmetic.CN.I_in\[29\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7322__S _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_506 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_517 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_528 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_539 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_87_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4847__I0 mod.Data_Mem.F_M.MRAM\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6461__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__I3 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6960__I _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7261__I1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4775__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5972__A1 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5576__I _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5724__A1 _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7791__I _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8539__D _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8130__RN net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout277_I net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4463__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5820_ _2347_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4215__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5751_ _1944_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4766__A2 mod.Arithmetic.ACTI.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4390__I _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4702_ _0661_ mod.Arithmetic.CN.I_in\[70\] _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8470_ _0566_ net237 mod.Data_Mem.F_M.MRAM\[796\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5682_ _2084_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7421_ mod.Data_Mem.F_M.MRAM\[776\]\[3\] _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8197__RN net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5715__A1 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4633_ mod.Arithmetic.CN.I_in\[37\] _1215_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7352_ _3649_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5191__A2 mod.Data_Mem.F_M.MRAM\[769\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4564_ _1111_ _1120_ _1234_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6303_ _2698_ _1967_ _2870_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7283_ _3232_ _3332_ _3604_ _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4495_ _1067_ _1072_ _1054_ _1056_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6110__I _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout92_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6234_ _2156_ _1842_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6140__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _2774_ _1685_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8509__572 net572 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ _1692_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5326__S0 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6096_ _2701_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8121__RN net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7491__I1 mod.Data_Mem.F_M.MRAM\[781\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5047_ _1711_ mod.Data_Mem.F_M.MRAM\[771\]\[1\] _1714_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4454__A1 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6780__I _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6998_ _3395_ mod.Data_Mem.F_M.MRAM\[17\]\[2\] _3435_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5954__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5949_ mod.Data_Mem.F_M.MRAM\[18\]\[5\] mod.Data_Mem.F_M.MRAM\[19\]\[5\] _2427_ _2569_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5396__I _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8337__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5706__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7619_ _3802_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5309__I1 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7116__I _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6131__A1 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6131__B2 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6682__A2 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7631__A1 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__A2 mod.Data_Mem.F_M.MRAM\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7482__I1 mod.Data_Mem.F_M.MRAM\[780\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8112__RN net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6690__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__A1 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5245__I0 mod.Data_Mem.F_M.MRAM\[771\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4748__A2 _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4280_ _0873_ _0650_ _0813_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_67_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4684__A1 mod.Arithmetic.CN.I_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8103__RN net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6425__A2 mod.Data_Mem.F_M.MRAM\[780\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7970_ _0196_ net79 mod.Data_Mem.F_M.MRAM\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7473__I1 mod.Data_Mem.F_M.MRAM\[780\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__A1 _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4436__B2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6921_ _3373_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7225__I1 mod.Data_Mem.F_M.MRAM\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _3348_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6189__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5210__S _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout18 net22 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5803_ _1835_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout29 net31 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_6783_ mod.Data_Mem.F_M.MRAM\[799\]\[1\] _3303_ _3300_ _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3995_ _0669_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6105__I _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8522_ _0026_ net340 mod.Data_Mem.F_M.out_data\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5734_ _2058_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8453_ _0549_ net315 mod.Data_Mem.F_M.MRAM\[794\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ _2264_ _2126_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7137__S _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4988__C _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _3675_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ _1205_ _1219_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8384_ _0480_ net180 mod.Data_Mem.F_M.MRAM\[785\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5596_ _2220_ _2228_ _2232_ _2218_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7335_ _3639_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6976__S _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4547_ _1207_ _1213_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7266_ _3595_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7161__I0 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _1044_ _1045_ _1143_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_89_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6217_ mod.Data_Mem.F_M.MRAM\[1\]\[3\] mod.Data_Mem.F_M.MRAM\[2\]\[3\] mod.Data_Mem.F_M.MRAM\[3\]\[3\]
+ mod.Data_Mem.F_M.MRAM\[4\]\[3\] _2632_ _2440_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_89_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7197_ _3555_ _3550_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _2757_ _2762_ _2763_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ _2695_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5155__A2 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7877__CLK net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__B _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6104__A1 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 mod.Arithmetic.CN.I_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4418__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4933__I _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5218__I0 _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5918__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__I0 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout142_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5764__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5450_ _1916_ _1495_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6343__A1 _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4401_ _1053_ _1057_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_126_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5381_ mod.Data_Mem.F_M.MRAM\[787\]\[7\] _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7120_ _3508_ mod.Data_Mem.F_M.MRAM\[3\]\[5\] _3506_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4332_ _0671_ _0848_ _0919_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__7143__I0 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout208 net212 net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7051_ _3472_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout219 net220 net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4263_ _0864_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8032__CLK net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6002_ _2406_ _2620_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5854__C2 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4194_ _0623_ _0656_ _0824_ _0839_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_80_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout55_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7953_ _0179_ net202 mod.Data_Mem.F_M.MRAM\[769\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6544__B _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5082__A1 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _3377_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7884_ _0110_ net376 mod.Data_Mem.F_M.MRAM\[26\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6835_ _3339_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ mod.Data_Mem.F_M.MRAM\[8\]\[6\] _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5385__A2 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3978_ _0635_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4999__B _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5717_ _2311_ _2152_ _2341_ _2342_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8505_ _0009_ net335 mod.Data_Mem.F_M.out_data\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6709__I0 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6697_ _3247_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5674__I _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8436_ _0532_ net155 mod.Data_Mem.F_M.MRAM\[792\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6334__A1 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5648_ _2063_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5137__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8367_ _0463_ net221 mod.Data_Mem.F_M.MRAM\[782\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5579_ mod.Data_Mem.F_M.MRAM\[797\]\[3\] _2176_ _2189_ mod.Data_Mem.F_M.MRAM\[796\]\[3\]
+ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7318_ _3555_ _3623_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7134__I0 _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8298_ _0394_ net196 mod.Data_Mem.F_M.MRAM\[773\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _3586_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6438__C _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6454__B _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4753__I mod.Arithmetic.CN.I_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5584__I _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6325__A1 mod.Data_Mem.F_M.MRAM\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6325__B2 mod.Data_Mem.F_M.MRAM\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7505__S _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__B1 mod.Data_Mem.F_M.MRAM\[791\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7825__A1 _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4928__I _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5151__I2 mod.Data_Mem.F_M.MRAM\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7240__S _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7053__A2 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6364__B _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout357_I net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A4 mod.Arithmetic.CN.I_in\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ _1507_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4811__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6939__I0 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4881_ _1536_ _1549_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6620_ _3200_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6564__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6564__B2 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _2338_ mod.Data_Mem.F_M.MRAM\[0\]\[7\] _2101_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5502_ _1791_ mod.Data_Mem.F_M.MRAM\[31\]\[6\] _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6316__A1 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6482_ _2133_ mod.Data_Mem.F_M.MRAM\[781\]\[3\] _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8221_ _0322_ net311 mod.Data_Mem.F_M.MRAM\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5433_ _2084_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8152_ mod.Data_Mem.F_M.out_data\[62\] net61 net362 mod.Arithmetic.CN.I_in\[62\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5364_ mod.Data_Mem.F_M.MRAM\[31\]\[7\] _1914_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7103_ _3498_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4315_ _0979_ _0987_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8083_ _0283_ net304 mod.Data_Mem.F_M.MRAM\[23\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5295_ mod.Data_Mem.F_M.MRAM\[771\]\[5\] mod.Data_Mem.F_M.MRAM\[770\]\[5\] _1874_
+ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5827__B1 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5827__C2 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7034_ _3461_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4246_ _0914_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6095__A3 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4177_ _0827_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5055__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7936_ _0162_ net341 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A1 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7867_ _0093_ net371 mod.Data_Mem.F_M.MRAM\[11\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6818_ mod.Data_Mem.F_M.MRAM\[789\]\[4\] _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7798_ _3897_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6749_ _3281_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8078__CLK net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4318__B1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8419_ _0515_ net138 mod.Data_Mem.F_M.MRAM\[790\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5353__B _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5133__I2 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__A1 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6963__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6184__B _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5046__A1 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6243__B1 _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__A2 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A1 _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6546__B2 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7594__I0 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4557__B1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4021__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout105_I net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4100_ _0753_ _0771_ _0775_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ _1517_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5285__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4031_ mod.Arithmetic.CN.I_in\[23\] _0683_ _0700_ _0706_ _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_84_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5982_ _2073_ _2601_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7721_ _3854_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4933_ _1601_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7652_ mod.Data_Mem.F_M.MRAM\[790\]\[2\] _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6537__A1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ mod.Data_Mem.F_M.src\[4\] _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6603_ mod.Data_Mem.F_M.MRAM\[11\]\[5\] _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7583_ _3780_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout18_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4795_ _1304_ _1320_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6534_ _3135_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5157__C _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5760__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _3065_ _3069_ _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8204_ _0305_ net296 mod.Data_Mem.F_M.MRAM\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5416_ _2073_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6396_ _2381_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8135_ mod.Data_Mem.F_M.out_data\[45\] net47 net279 mod.Arithmetic.CN.I_in\[45\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5347_ _1923_ mod.Data_Mem.F_M.MRAM\[786\]\[6\] _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8066_ _0275_ net186 mod.Data_Mem.F_M.MRAM\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5278_ _1830_ _1941_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5276__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7017_ _3239_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4229_ _0902_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__A1 _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7919_ _0145_ net201 mod.Data_Mem.F_M.MRAM\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6528__A1 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6379__I1 mod.Data_Mem.F_M.MRAM\[791\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7576__I0 _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7119__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5200__A1 mod.Data_Mem.F_M.MRAM\[799\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6023__I _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6000__I0 mod.Data_Mem.F_M.MRAM\[770\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5503__A2 mod.Data_Mem.F_M.MRAM\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5267__B2 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout380 net381 net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__S _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5362__S1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout391 net392 net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5019__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__A2 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A2 mod.Arithmetic.ACTI.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4941__I _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8560__D _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7567__I0 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5990__A2 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout222_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ _1061_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6250_ _2523_ _2840_ _2860_ _2863_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ _1758_ mod.Data_Mem.F_M.MRAM\[15\]\[3\] mod.Data_Mem.F_M.MRAM\[31\]\[3\] _1724_
+ _1675_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4388__I _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6181_ _1589_ _2795_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5132_ _1796_ mod.Data_Mem.F_M.MRAM\[785\]\[2\] _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _1730_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6309__S _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _0637_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_37_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5012__I _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5965_ _2499_ _2583_ _2584_ _2555_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5430__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__I1 mod.Data_Mem.F_M.MRAM\[786\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7704_ mod.Data_Mem.F_M.MRAM\[793\]\[4\] _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4916_ _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5896_ mod.Data_Mem.F_M.MRAM\[16\]\[3\] mod.Data_Mem.F_M.MRAM\[17\]\[3\] _2516_ _2518_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5168__B _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3992__A1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7635_ _3811_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4847_ mod.Data_Mem.F_M.MRAM\[19\]\[0\] mod.Data_Mem.F_M.MRAM\[18\]\[0\] _1515_ _1516_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7566_ _3769_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4778_ _1310_ _1318_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6778__I _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6517_ _3030_ _2323_ _3023_ _2569_ _2572_ _3022_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_106_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7497_ _3725_ mod.Data_Mem.F_M.MRAM\[781\]\[4\] _3726_ _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _2689_ mod.Data_Mem.F_M.MRAM\[780\]\[2\] _2375_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8116__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5497__A1 _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4298__I _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6379_ mod.Data_Mem.F_M.MRAM\[789\]\[7\] mod.Data_Mem.F_M.MRAM\[791\]\[7\] mod.Data_Mem.F_M.MRAM\[790\]\[7\]
+ mod.Data_Mem.F_M.MRAM\[788\]\[7\] _2167_ _2376_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_103_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__S _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8118_ mod.Data_Mem.F_M.out_data\[28\] net41 net274 mod.Arithmetic.CN.I_in\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_507 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_518 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_8049_ _0258_ net209 mod.Data_Mem.F_M.MRAM\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_529 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__I1 mod.Data_Mem.F_M.MRAM\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__I0 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4224__A2 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5972__A2 mod.Data_Mem.F_M.MRAM\[772\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3983__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5592__I _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7513__S _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4160__A1 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8555__D _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7312__I _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5660__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4463__A2 mod.Arithmetic.CN.I_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4215__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _2374_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4701_ _1370_ _1248_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5681_ _2309_ mod.Data_Mem.F_M.MRAM\[29\]\[4\] _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7420_ _3683_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4632_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__A2 mod.Data_Mem.F_M.MRAM\[797\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5716__B _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4563_ _1111_ _1120_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7351_ mod.Data_Mem.F_M.MRAM\[772\]\[0\] _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6302_ _2868_ _1966_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7282_ _3297_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4494_ _1052_ _1074_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5479__A1 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6233_ _1936_ _1848_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__I _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _1608_ _1691_ _2733_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _1598_ _1779_ _1781_ _1509_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6039__S _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6095_ _2704_ _2682_ _2711_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5326__S1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _1712_ _1713_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5651__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__A2 mod.Arithmetic.ACTI.x\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6997_ _3437_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5403__A1 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _2523_ _2545_ _2568_ _2407_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_34_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5954__A2 mod.Data_Mem.F_M.MRAM\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ _2296_ mod.Data_Mem.F_M.MRAM\[771\]\[3\] _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7618_ _3749_ mod.Data_Mem.F_M.MRAM\[787\]\[2\] _3801_ _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5706__A2 mod.Data_Mem.F_M.MRAM\[796\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7549_ _3232_ _3298_ _3758_ _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5309__I2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6131__A2 mod.Data_Mem.F_M.MRAM\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4142__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4693__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7631__A2 _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5642__A1 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5587__I _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5245__I1 mod.Data_Mem.F_M.MRAM\[770\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A2 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6412__S _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5253__S0 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8431__CLK net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4133__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8581__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout387_I net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4436__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6881__I mod.Data_Mem.F_M.MRAM\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6920_ _3227_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6851_ mod.Data_Mem.F_M.MRAM\[779\]\[1\] _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6189__A2 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5802_ _2107_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout19 net22 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_90_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6782_ _3302_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3994_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8521_ _0025_ net332 mod.Data_Mem.F_M.out_data\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4995__I0 mod.Data_Mem.F_M.MRAM\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ mod.Data_Mem.F_M.MRAM\[18\]\[0\] mod.Data_Mem.F_M.MRAM\[19\]\[0\] _2297_ _2358_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8452_ _0548_ net375 mod.Data_Mem.F_M.MRAM\[794\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5664_ _2068_ _2117_ _2288_ _2294_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7403_ mod.Data_Mem.F_M.MRAM\[775\]\[2\] _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4747__I0 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4615_ _1284_ _1195_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8383_ _0479_ net117 mod.Data_Mem.F_M.MRAM\[784\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5595_ mod.Data_Mem.F_M.MRAM\[797\]\[4\] _2214_ _1750_ mod.Data_Mem.F_M.MRAM\[796\]\[4\]
+ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7217__I _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6361__A2 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7334_ _3638_ mod.Data_Mem.F_M.MRAM\[771\]\[1\] _3636_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4546_ _1214_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7265_ mod.Data_Mem.F_M.MRAM\[5\]\[0\] _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4477_ _0731_ _0722_ _0820_ _0972_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_104_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7161__I1 mod.Data_Mem.F_M.MRAM\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6216_ _2828_ _2829_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7196_ _3308_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5872__A1 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6147_ _2178_ _1659_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6078_ _2202_ _2194_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ _1693_ mod.Data_Mem.F_M.MRAM\[791\]\[1\] _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8304__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7127__I _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5560__B1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5870__I _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8097__RN net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4418__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5218__I1 _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__I1 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__A1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7238__S _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout135_I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6343__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4400_ _1067_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout302_I net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ _1703_ _2041_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5551__B1 mod.Data_Mem.F_M.MRAM\[798\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4331_ _0912_ _0919_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7143__I1 mod.Data_Mem.F_M.MRAM\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5154__I0 mod.Data_Mem.F_M.MRAM\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7050_ _3456_ mod.Data_Mem.F_M.MRAM\[1\]\[4\] _3469_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout209 net211 net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4262_ _0867_ _0936_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6001_ _2102_ _2619_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5854__B2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4193_ _0816_ _0821_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__A1 mod.Data_Mem.F_M.MRAM\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__B2 mod.Data_Mem.F_M.MRAM\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7952_ _0178_ net201 mod.Data_Mem.F_M.MRAM\[769\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5082__A2 _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6903_ _3228_ mod.Data_Mem.F_M.MRAM\[13\]\[0\] _3376_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout48_I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7883_ _0109_ net384 mod.Data_Mem.F_M.MRAM\[26\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6116__I _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6834_ _3240_ mod.Data_Mem.F_M.MRAM\[769\]\[1\] _3337_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8477__CLK net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _3289_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6582__A2 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3977_ _0619_ mod.Arithmetic.CN.I_in\[32\] _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7148__S _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8504_ _0008_ net349 mod.Data_Mem.F_M.out_data\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6052__S _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ _2157_ mod.Data_Mem.F_M.MRAM\[796\]\[7\] _2210_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ _3246_ mod.Data_Mem.F_M.MRAM\[28\]\[3\] _3237_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6709__I1 mod.Data_Mem.F_M.MRAM\[28\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5176__B _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8435_ _0531_ net377 mod.Data_Mem.F_M.MRAM\[792\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6987__S _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5647_ _2278_ mod.Data_Mem.F_M.MRAM\[29\]\[1\] _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5891__S _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6334__A2 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4345__A1 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8366_ _0462_ net221 mod.Data_Mem.F_M.MRAM\[782\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5542__B1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _2214_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6786__I _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7317_ _1770_ _3626_ _3628_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4529_ _1198_ _1199_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7134__I1 mod.Data_Mem.F_M.MRAM\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8297_ _0393_ net185 mod.Data_Mem.F_M.MRAM\[773\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6098__A1 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7248_ mod.Data_Mem.F_M.MRAM\[31\]\[0\] _3293_ _3585_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5845__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4648__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7179_ mod.Data_Mem.F_M.MRAM\[22\]\[4\] _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7598__A1 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8079__RN net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6454__C _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5865__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4336__A1 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6089__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__B2 _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5836__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5151__I3 mod.Data_Mem.F_M.MRAM\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8563__D _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5041__S _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6261__A1 _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout252_I net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ mod.Data_Mem.F_M.MRAM\[3\]\[0\] _1539_ _1540_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6939__I1 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5775__I _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__A2 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6550_ _2722_ mod.Data_Mem.F_M.MRAM\[1\]\[7\] _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5501_ _2081_ _2140_ _2144_ _2102_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6481_ _2635_ _3086_ _1623_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8220_ _0321_ net311 mod.Data_Mem.F_M.MRAM\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4327__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5375__I0 mod.Data_Mem.F_M.MRAM\[773\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5432_ _1493_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5363_ _1888_ _2024_ _1884_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8151_ mod.Data_Mem.F_M.out_data\[61\] net61 net361 mod.Arithmetic.CN.I_in\[61\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_114_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5216__S _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7102_ mod.Data_Mem.F_M.MRAM\[23\]\[6\] _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _0979_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5294_ _1954_ _1955_ _1957_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8082_ _0282_ net141 mod.Data_Mem.F_M.MRAM\[23\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5827__B2 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7033_ _3460_ mod.Data_Mem.F_M.MRAM\[18\]\[6\] _3457_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4245_ _0912_ _0915_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_68_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4176_ _0829_ _0840_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_67_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7935_ _0161_ net339 mod.Data_Mem.F_M.MRAM\[799\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7866_ _0092_ net167 mod.Data_Mem.F_M.MRAM\[11\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _3327_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7797_ _3319_ mod.Data_Mem.F_M.MRAM\[798\]\[6\] _3894_ _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4566__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ _3253_ mod.Data_Mem.F_M.MRAM\[0\]\[5\] _3279_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4566__B2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6679_ mod.DMen_reg2 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4318__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8418_ _0514_ net188 mod.Data_Mem.F_M.MRAM\[790\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5366__I0 mod.Data_Mem.F_M.MRAM\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4318__B2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8349_ _0445_ net230 mod.Data_Mem.F_M.MRAM\[780\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7405__I mod.Data_Mem.F_M.MRAM\[775\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5133__I3 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__A2 _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__B _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__I0 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6546__A2 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4557__A1 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4004__I mod.Arithmetic.CN.I_in\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4309__A1 _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5506__B1 _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8172__CLK net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8558__D _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4939__I _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5263__C _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5809__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4875__S _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4030_ _0702_ mod.Arithmetic.I_out\[78\] _0703_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6234__A1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _1633_ _2593_ _2594_ _2102_ _2557_ _2600_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_80_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7720_ mod.Data_Mem.F_M.MRAM\[794\]\[4\] _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ _1524_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7651_ _3819_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ _1497_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6537__A2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6602_ _3191_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7582_ _3778_ mod.Data_Mem.F_M.MRAM\[785\]\[4\] _3779_ _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4794_ _1423_ _1332_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6533_ _2252_ mod.Data_Mem.F_M.MRAM\[0\]\[6\] _2100_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7337__I1 mod.Data_Mem.F_M.MRAM\[771\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _2827_ _3070_ _2080_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8203_ _0304_ net297 mod.Data_Mem.F_M.MRAM\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5415_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4849__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6395_ _2419_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6269__C _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8134_ mod.Data_Mem.F_M.out_data\[44\] net44 net255 mod.Arithmetic.CN.I_in\[44\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5346_ mod.Data_Mem.F_M.MRAM\[787\]\[6\] _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8065_ _0274_ net148 mod.Data_Mem.F_M.MRAM\[21\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5277_ mod.Data_Mem.F_M.MRAM\[791\]\[5\] mod.Data_Mem.F_M.MRAM\[790\]\[5\] _1512_
+ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7161__S _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5276__A2 mod.Data_Mem.F_M.MRAM\[789\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6473__A1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7016_ _3449_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4228_ _0892_ _0901_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4159_ _0834_ mod.Arithmetic.CN.I_in\[41\] _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6225__A1 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7918_ _0144_ net207 mod.Data_Mem.F_M.MRAM\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4787__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7849_ mod.Data_Mem.F_M.MRAM\[9\]\[3\] _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6528__A2 _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4539__A1 mod.Arithmetic.CN.I_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8195__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5200__A2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5339__I0 mod.Data_Mem.F_M.MRAM\[773\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6000__I1 mod.Data_Mem.F_M.MRAM\[771\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6839__I0 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6464__A1 _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout370 net374 net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout381 net389 net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout392 net393 net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__A2 _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__I1 mod.Data_Mem.F_M.MRAM\[784\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout215_I net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__I _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5200_ mod.Data_Mem.F_M.MRAM\[799\]\[3\] _1635_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4702__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6180_ _2064_ mod.Data_Mem.F_M.MRAM\[14\]\[2\] mod.Data_Mem.F_M.MRAM\[15\]\[2\] _2095_
+ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5131_ _1792_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6455__A1 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5889__S0 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5062_ _1632_ _1677_ _1729_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4013_ mod.Arithmetic.CN.I_in\[17\] _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8068__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4769__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ mod.Data_Mem.F_M.MRAM\[14\]\[5\] mod.Data_Mem.F_M.MRAM\[15\]\[5\] _2516_ _2584_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7007__I0 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7703_ _3845_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout30_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5430__A2 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4915_ _1583_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5895_ mod.Data_Mem.F_M.MRAM\[14\]\[3\] mod.Data_Mem.F_M.MRAM\[15\]\[3\] _2516_ _2517_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7634_ mod.Data_Mem.F_M.MRAM\[788\]\[1\] _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5718__B1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4846_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3992__A2 mod.Arithmetic.CN.I_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7905__CLK net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5194__A1 _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ _3729_ mod.Data_Mem.F_M.MRAM\[784\]\[6\] _3759_ _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _1298_ _1445_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6516_ _3114_ _3116_ _3119_ _3013_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7496_ _3719_ _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4579__I mod.Arithmetic.CN.I_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6447_ _3016_ mod.Data_Mem.F_M.MRAM\[781\]\[2\] _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5497__A2 mod.Data_Mem.F_M.MRAM\[30\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6378_ _2883_ _2984_ _2987_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8117_ mod.Data_Mem.F_M.out_data\[27\] net46 net329 mod.Arithmetic.CN.I_in\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5329_ mod.Data_Mem.F_M.MRAM\[23\]\[6\] mod.Data_Mem.F_M.MRAM\[22\]\[6\] _1890_ _1992_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6446__A1 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_508 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_8048_ _0257_ net207 mod.Data_Mem.F_M.MRAM\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_519 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__I1 mod.Data_Mem.F_M.MRAM\[798\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3983__A2 mod.Arithmetic.CN.I_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5732__I0 mod.Data_Mem.F_M.MRAM\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4160__A2 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5314__S _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5113__I _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5660__A2 mod.Data_Mem.F_M.MRAM\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__I1 mod.Data_Mem.F_M.MRAM\[798\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8571__D _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5948__B1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout165_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout332_I net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4700_ _1243_ _1247_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5680_ _1693_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _1169_ _1183_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5176__A1 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7350_ _3648_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4923__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4562_ _1225_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _2864_ _2913_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7281_ _3292_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4493_ _1049_ _1163_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5479__A2 _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6232_ _2841_ _2843_ _2732_ _2845_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6163_ _1920_ _1697_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7476__I0 _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5114_ mod.Data_Mem.F_M.MRAM\[783\]\[2\] _1780_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout78_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6094_ _2189_ _2706_ _2707_ _2710_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5045_ mod.Data_Mem.F_M.MRAM\[770\]\[1\] _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5651__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4454__A3 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _3393_ mod.Data_Mem.F_M.MRAM\[17\]\[1\] _3435_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5403__A2 _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5947_ _2520_ _2556_ _2567_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5878_ _1791_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7617_ _3797_ _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6789__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4829_ _1494_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7548_ _3420_ _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7479_ _3715_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5309__I3 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8233__CLK net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4142__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3941__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6419__A1 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8383__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5642__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5868__I _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5158__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6355__B1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5253__S1 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7524__S _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4133__A2 mod.Arithmetic.CN.I_in\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout282_I net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _3347_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5801_ _1535_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8106__CLK net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6781_ net4 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3993_ _0632_ mod.Arithmetic.ACTI.x\[0\] _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8520_ _0024_ net350 mod.Data_Mem.F_M.out_data\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5732_ mod.Data_Mem.F_M.MRAM\[4\]\[0\] mod.Data_Mem.F_M.MRAM\[5\]\[0\] mod.Data_Mem.F_M.MRAM\[20\]\[0\]
+ mod.Data_Mem.F_M.MRAM\[21\]\[0\] _1717_ _1757_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4995__I1 mod.Data_Mem.F_M.MRAM\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8451_ _0547_ net377 mod.Data_Mem.F_M.MRAM\[794\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5663_ _2062_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7402_ _3674_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _1165_ _1187_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8382_ _0478_ net116 mod.Data_Mem.F_M.MRAM\[784\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4747__I1 mod.Arithmetic.CN.I_in\[70\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5594_ _1708_ _2230_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7333_ _3302_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4545_ _1215_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7264_ _3594_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _1031_ _1032_ _1034_ _1148_ mod.P3.Res\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_89_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6215_ _2558_ _2510_ mod.Data_Mem.F_M.MRAM\[20\]\[3\] _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5321__A1 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _3554_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__A2 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6146_ _1752_ _1663_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6077_ _2076_ _1498_ _2161_ _1633_ _2693_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5624__A2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5028_ _1695_ mod.Data_Mem.F_M.MRAM\[790\]\[1\] _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__A1 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _3426_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7609__S _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3936__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4033__S _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5560__A1 mod.Data_Mem.F_M.MRAM\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5560__B2 mod.Data_Mem.F_M.MRAM\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6468__B _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6982__I _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8129__CLK net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5218__I2 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6040__A2 mod.Data_Mem.F_M.MRAM\[21\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4007__I mod.Arithmetic.CN.I_in\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6328__B1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5039__S _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout128_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__A1 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__B2 _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__S _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4330_ _0921_ _0926_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5154__I1 mod.Data_Mem.F_M.MRAM\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4261_ _0868_ _0888_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6500__B1 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ mod.Data_Mem.F_M.MRAM\[770\]\[6\] mod.Data_Mem.F_M.MRAM\[771\]\[6\] _2271_
+ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5854__A2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4192_ _0865_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input2_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7951_ _0177_ net187 mod.Data_Mem.F_M.MRAM\[769\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _3375_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7882_ _0108_ net155 mod.Data_Mem.F_M.MRAM\[26\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4290__A1 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7603__I0 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _3338_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ mod.Data_Mem.F_M.MRAM\[8\]\[5\] _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ _0631_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8503_ _0007_ net246 mod.Data_Mem.F_M.out_data\[79\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5715_ _2278_ mod.Data_Mem.F_M.MRAM\[797\]\[7\] _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6695_ _3245_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7228__I _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8434_ _0530_ net323 mod.Data_Mem.F_M.MRAM\[792\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5646_ _2094_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8365_ _0461_ net229 mod.Data_Mem.F_M.MRAM\[782\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4345__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5542__A1 mod.Data_Mem.F_M.MRAM\[797\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5577_ _1783_ mod.Data_Mem.F_M.MRAM\[799\]\[3\] mod.Data_Mem.F_M.MRAM\[798\]\[3\]
+ _2084_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7316_ _3612_ _3623_ _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4528_ _1108_ _1140_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8296_ _0392_ net151 mod.Data_Mem.F_M.MRAM\[773\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7295__A1 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6098__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7247_ _3584_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_78_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4459_ _1125_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7178_ _3544_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6129_ _1537_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7598__A2 _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4281__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5211__I _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__B1 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__S _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__I0 mod.Data_Mem.F_M.MRAM\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8571__CLK net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4336__A2 mod.Arithmetic.ACTI.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5384__I1 mod.Data_Mem.F_M.MRAM\[784\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__I _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A2 mod.Data_Mem.F_M.MRAM\[790\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5836__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5322__S _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6261__A2 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6549__B1 _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout245_I net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ _2141_ _2143_ _2067_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _3084_ _1855_ _3085_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6887__I mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5431_ _2057_ _0010_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5375__I1 mod.Data_Mem.F_M.MRAM\[772\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4327__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5791__I _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8150_ mod.Data_Mem.F_M.out_data\[60\] net62 net363 mod.Arithmetic.CN.I_in\[60\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5362_ _2020_ _2021_ _2022_ _2023_ _1698_ _1664_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ _3497_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ _0982_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8081_ _0281_ net140 mod.Data_Mem.F_M.MRAM\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5293_ _1956_ mod.Data_Mem.F_M.MRAM\[768\]\[5\] _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5827__A2 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7032_ _3255_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _0916_ _0918_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4175_ _0841_ _0843_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_67_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout60_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7934_ _0160_ net332 mod.Data_Mem.F_M.MRAM\[799\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7865_ _0091_ net166 mod.Data_Mem.F_M.MRAM\[11\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4870__I _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ mod.Data_Mem.F_M.MRAM\[789\]\[3\] _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7796_ _3896_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6998__S _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6747_ _3280_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4566__A2 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3959_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7992__RN net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6678_ _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5629_ _1494_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8417_ _0513_ net150 mod.Data_Mem.F_M.MRAM\[790\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5366__I1 mod.Data_Mem.F_M.MRAM\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8348_ _0444_ net230 mod.Data_Mem.F_M.MRAM\[780\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8279_ _0375_ net121 mod.Data_Mem.F_M.MRAM\[770\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4110__I mod.Arithmetic.ACTI.x\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6243__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6481__B _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5876__I _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__I1 mod.Data_Mem.F_M.MRAM\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5754__A1 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6701__S _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7983__RN net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5506__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4309__A2 mod.Arithmetic.CN.I_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5506__B2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4020__I mod.Arithmetic.CN.I_in\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8574__D _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6482__A2 mod.Data_Mem.F_M.MRAM\[781\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4955__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout195_I net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5980_ _2387_ _2140_ _2390_ _2596_ _2599_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_80_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _1599_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5786__I _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7650_ mod.Data_Mem.F_M.MRAM\[790\]\[1\] _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4862_ mod.Data_Mem.F_M.MRAM\[22\]\[0\] _1513_ _1516_ _1520_ _1526_ _1530_ _1531_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_60_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6537__A3 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6601_ mod.Data_Mem.F_M.MRAM\[11\]\[4\] _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7581_ _3772_ _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5745__A1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4793_ _1422_ _1462_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6532_ _2289_ mod.Data_Mem.F_M.MRAM\[1\]\[6\] _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _3047_ _2293_ _3008_ _2476_ _2480_ _2484_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_8202_ _0087_ net12 net115 mod.I_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5414_ _1673_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6410__I _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6170__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6394_ _2090_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8133_ mod.Data_Mem.F_M.out_data\[43\] net47 net279 mod.Arithmetic.CN.I_in\[43\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _1732_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5026__I _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8064_ _0273_ net147 mod.Data_Mem.F_M.MRAM\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5276_ _1937_ mod.Data_Mem.F_M.MRAM\[789\]\[5\] _1939_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7015_ _3445_ mod.Data_Mem.F_M.MRAM\[18\]\[0\] _3448_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4227_ _0892_ _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6285__C _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _0618_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4089_ _0742_ _0748_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7984__CLK net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7917_ _0143_ net174 mod.Data_Mem.F_M.MRAM\[10\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7848_ _3926_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6379__I3 mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4539__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7779_ _3886_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4105__I _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5339__I1 mod.Data_Mem.F_M.MRAM\[772\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3944__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4041__S _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6161__A1 _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6839__I1 mod.Data_Mem.F_M.MRAM\[769\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout360 net366 net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout371 net373 net371 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xfanout382 net385 net382 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout393 net1 net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6216__A2 _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout110_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout208_I net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4702__A2 mod.Arithmetic.CN.I_in\[70\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ mod.Data_Mem.F_M.MRAM\[784\]\[2\] _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5889__S1 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8133__RN net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5061_ _1701_ _1726_ _1728_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4012_ mod.Arithmetic.I_out\[74\] _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_96_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6207__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4218__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5963_ mod.Data_Mem.F_M.MRAM\[2\]\[5\] mod.Data_Mem.F_M.MRAM\[3\]\[5\] _2582_ _2583_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5966__A1 _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4769__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4634__B _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7007__I1 mod.Data_Mem.F_M.MRAM\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7702_ mod.Data_Mem.F_M.MRAM\[793\]\[3\] _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4914_ _1541_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5894_ _1944_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA_fanout23_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5718__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4845_ _1510_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7633_ _3810_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5718__B2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6341__S _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7564_ _3768_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4776_ _1301_ _1322_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6515_ _3059_ _2583_ _2584_ _3019_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7495_ _3311_ _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6143__A1 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6446_ _3002_ _3052_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7191__I0 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6377_ _2727_ _2985_ _2986_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8116_ mod.Data_Mem.F_M.out_data\[26\] net52 net334 mod.Arithmetic.CN.I_in\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5328_ mod.Data_Mem.F_M.MRAM\[31\]\[6\] _1886_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8047_ _0256_ net207 mod.Data_Mem.F_M.MRAM\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8124__RN net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_509 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_5259_ _1923_ mod.Data_Mem.F_M.MRAM\[786\]\[4\] _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8012__CLK net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4209__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8162__CLK net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3939__I _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7347__S _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6134__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5732__I1 mod.Data_Mem.F_M.MRAM\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4696__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8115__RN net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout190 net194 net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_94_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8505__CLK net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5330__S _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A1 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6996__I0 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout158_I net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__I0 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7257__S _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout325_I net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4630_ _1166_ _1299_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6373__A1 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5176__A2 mod.Data_Mem.F_M.MRAM\[775\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4561_ _1227_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4923__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _2866_ _2899_ _2912_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7280_ _3602_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6125__A1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4492_ _1075_ _1076_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6231_ _2156_ _1826_ _2771_ _2844_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _2771_ _2773_ _2777_ _2685_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4151__A3 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6428__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _1597_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7476__I1 mod.Data_Mem.F_M.MRAM\[780\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8106__RN net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _2709_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5044_ _1542_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5240__S _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6563__C _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5939__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6987__I0 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _3436_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _2557_ _2561_ _2564_ _2566_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6739__I0 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5877_ _2498_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4828_ _1495_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7616_ _3800_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6364__A1 _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7547_ _3757_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4759_ _1418_ _1420_ _1428_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_111_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7478_ _3645_ mod.Data_Mem.F_M.MRAM\[780\]\[5\] _3713_ _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6429_ _2550_ _2429_ _3036_ _2498_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4602__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5884__I _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6355__A1 mod.Data_Mem.F_M.MRAM\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6355__B2 mod.Data_Mem.F_M.MRAM\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6107__A1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5325__S _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4669__A1 mod.Arithmetic.CN.I_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5124__I _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4963__I _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8582__D _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout275_I net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5800_ _2413_ _2423_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6780_ _3301_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3992_ _0668_ mod.Arithmetic.CN.I_in\[64\] _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5731_ _2110_ _2348_ _2350_ _2352_ _2354_ _2355_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5794__I _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8450_ _0546_ net167 mod.Data_Mem.F_M.MRAM\[794\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6346__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5662_ _2290_ _2291_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7401_ mod.Data_Mem.F_M.MRAM\[775\]\[1\] _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4613_ _1165_ _1187_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8381_ _0477_ net110 mod.Data_Mem.F_M.MRAM\[784\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5593_ _2229_ mod.Data_Mem.F_M.MRAM\[799\]\[4\] mod.Data_Mem.F_M.MRAM\[798\]\[4\]
+ _1816_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7332_ _3637_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4544_ mod.Arithmetic.CN.I_in\[35\] _1091_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7263_ mod.Data_Mem.F_M.MRAM\[31\]\[7\] _3322_ _3590_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4475_ _1031_ _1146_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6214_ _2205_ _2212_ _2496_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout90_I net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7194_ _3529_ mod.Data_Mem.F_M.MRAM\[29\]\[2\] _3553_ _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5321__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _2744_ _2756_ _2760_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5034__I _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__B1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _2079_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4873__I _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _1694_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__B _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6978_ _3395_ mod.Data_Mem.F_M.MRAM\[16\]\[2\] _3423_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _2389_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8200__CLK net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6337__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8579_ _0595_ net218 mod.Instr_Mem.instruction\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5209__I _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7137__I0 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5560__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5848__B1 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4984__S _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5218__I3 _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5828__B _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6328__A1 mod.Data_Mem.F_M.MRAM\[781\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6328__B2 mod.Data_Mem.F_M.MRAM\[780\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5119__I _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7128__I0 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__A2 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__B1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4260_ _0891_ _0904_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6500__A1 _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6500__B2 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout392_I net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4191_ _0823_ _0853_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7300__I0 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7950_ _0176_ net187 mod.Data_Mem.F_M.MRAM\[769\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6901_ _3235_ _3371_ _3374_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7881_ _0107_ net321 mod.Data_Mem.F_M.MRAM\[26\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4290__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _3228_ mod.Data_Mem.F_M.MRAM\[769\]\[0\] _3337_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7603__I1 mod.Data_Mem.F_M.MRAM\[786\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8223__CLK net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6567__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _3288_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3975_ _0638_ _0651_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8502_ _0006_ net264 mod.Data_Mem.F_M.out_data\[78\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5714_ _2308_ _2150_ _2336_ _2339_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6319__A1 _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6694_ net6 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8433_ _0529_ net193 mod.Data_Mem.F_M.MRAM\[792\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5645_ _1494_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8364_ _0460_ net221 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5576_ _1554_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5542__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7315_ _1713_ _3626_ _3627_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4527_ _1108_ _1140_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4868__I _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8295_ _0391_ net83 mod.Data_Mem.F_M.MRAM\[772\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7295__A2 _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7246_ _3294_ _3464_ _3296_ _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4458_ _1126_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7177_ mod.Data_Mem.F_M.MRAM\[22\]\[3\] _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4389_ mod.Arithmetic.CN.I_in\[28\] _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6128_ _2684_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A1 mod.Data_Mem.F_M.MRAM\[783\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6059_ _2506_ mod.Data_Mem.F_M.MRAM\[782\]\[0\] mod.Data_Mem.F_M.MRAM\[783\]\[0\]
+ _2558_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_86_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A1 _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6558__B2 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3947__I _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4336__A3 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6993__I _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5830__C _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5402__I _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5844__I0 mod.Data_Mem.F_M.MRAM\[782\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6549__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout140_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout238_I net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7349__I0 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ _2074_ _2071_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5361_ mod.Data_Mem.F_M.MRAM\[7\]\[7\] mod.Data_Mem.F_M.MRAM\[6\]\[7\] _1890_ _2023_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7064__I mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4312_ _0984_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7100_ mod.Data_Mem.F_M.MRAM\[23\]\[5\] _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8080_ _0280_ net160 mod.Data_Mem.F_M.MRAM\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5292_ _1651_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7031_ _3459_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4243_ _0846_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_45_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__C _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4174_ _0666_ _0845_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_83_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout53_I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7933_ _0159_ net166 mod.Data_Mem.F_M.MRAM\[8\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5460__A1 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7864_ _0090_ net173 mod.Data_Mem.F_M.MRAM\[11\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _3326_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4015__A2 mod.Arithmetic.I_out\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7795_ _3806_ mod.Data_Mem.F_M.MRAM\[798\]\[5\] _3894_ _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6746_ _3249_ mod.Data_Mem.F_M.MRAM\[0\]\[4\] _3279_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3958_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5763__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6677_ mod.Data_Mem.F_M.dest\[1\] mod.Data_Mem.F_M.dest\[0\] _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8416_ _0512_ net149 mod.Data_Mem.F_M.MRAM\[790\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5628_ _1956_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8347_ _0443_ net254 mod.Data_Mem.F_M.MRAM\[780\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5559_ _1657_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8278_ _0374_ net121 mod.Data_Mem.F_M.MRAM\[770\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5279__A1 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _3523_ mod.Data_Mem.F_M.MRAM\[30\]\[0\] _3574_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__I0 mod.Data_Mem.F_M.MRAM\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5378__B _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5754__A2 mod.Data_Mem.F_M.MRAM\[769\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5506__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7612__I _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6228__I _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout188_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4245__A2 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _1523_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout355_I net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__A2 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6600_ _3190_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7580_ _3311_ _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4792_ _0702_ _1460_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5745__A2 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6898__I mod.Data_Mem.F_M.dest\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6531_ _2562_ mod.Data_Mem.F_M.MRAM\[13\]\[6\] _3115_ _3133_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6462_ _3067_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8201_ _0086_ net12 net114 mod.I_addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5413_ _2066_ _2068_ _2071_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6393_ _2617_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6170__A2 _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5344_ _1703_ _2006_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8132_ mod.Data_Mem.F_M.out_data\[42\] net46 net327 mod.Arithmetic.CN.I_in\[42\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8063_ _0272_ net163 mod.Data_Mem.F_M.MRAM\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5275_ _1921_ _1938_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7014_ _3447_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4226_ _0896_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6473__A3 _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4484__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5681__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4157_ _0831_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5042__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4088_ _0763_ _0764_ _0739_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7916_ _0142_ net172 mod.Data_Mem.F_M.MRAM\[10\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3995__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7847_ mod.Data_Mem.F_M.MRAM\[9\]\[2\] _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8519__566 net566 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7778_ _3782_ mod.Data_Mem.F_M.MRAM\[797\]\[6\] _3883_ _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5926__B _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ mod.Data_Mem.F_M.MRAM\[10\]\[7\] _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8091__CLK net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4172__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3960__I mod.Arithmetic.CN.I_in\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout350 net351 net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout361 net364 net361 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout372 net373 net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout383 net384 net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_93_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5975__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6511__I _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout103_I net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8584__CLK net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4966__I mod.Data_Mem.F_M.MRAM\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _1727_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4011_ mod.Arithmetic.CN.I_in\[18\] _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4466__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5663__A1 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4218__A2 mod.Arithmetic.CN.I_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _1512_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4634__C _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4769__A3 mod.Arithmetic.CN.I_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7701_ _3844_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3977__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4913_ _1581_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5893_ _2204_ _2514_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7632_ mod.Data_Mem.F_M.MRAM\[788\]\[0\] _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4844_ mod.Data_Mem.F_M.MRAM\[21\]\[0\] mod.Data_Mem.F_M.MRAM\[20\]\[0\] _1512_ _1513_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5718__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout16_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7563_ _3754_ mod.Data_Mem.F_M.MRAM\[784\]\[5\] _3760_ _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6391__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4775_ _1301_ _1322_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7517__I _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6514_ _2418_ _1968_ _2399_ _3117_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7494_ _3724_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6445_ _3030_ _2287_ _3004_ _2456_ _2459_ _3022_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__6143__A2 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7191__I1 mod.Data_Mem.F_M.MRAM\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4154__A1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6376_ _1638_ _2038_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8115_ mod.Data_Mem.F_M.out_data\[25\] net51 net337 mod.Arithmetic.CN.I_in\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_102_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5327_ _1872_ _1989_ _1884_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7951__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8046_ _0255_ net106 mod.Data_Mem.F_M.MRAM\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5258_ _1694_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5654__A1 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4209_ _0817_ _0721_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ mod.Data_Mem.F_M.MRAM\[768\]\[3\] _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8307__CLK net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4209__A2 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3968__A1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4768__I0 mod.Arithmetic.ACTI.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3955__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A1 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5893__A1 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout180 net181 net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout191 net194 net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5410__I _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6996__I1 mod.Data_Mem.F_M.MRAM\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6070__A1 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4620__A2 mod.Arithmetic.CN.I_in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6748__I1 mod.Data_Mem.F_M.MRAM\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6373__A2 _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout220_I net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__I _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4384__A1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4560_ _1228_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_fanout318_I net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4491_ _1075_ _1076_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_128_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4136__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6230_ _1740_ _1828_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6161_ _2702_ _2775_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7072__I mod.Data_Mem.F_M.MRAM\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5112_ _1566_ _1766_ _1773_ _1778_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _2708_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4439__A2 mod.Arithmetic.CN.I_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6684__I0 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4645__B _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6994_ _3386_ mod.Data_Mem.F_M.MRAM\[17\]\[0\] _3435_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5939__A2 mod.Data_Mem.F_M.MRAM\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6987__I1 mod.Data_Mem.F_M.MRAM\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6061__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _2562_ _1870_ _2069_ _2565_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4611__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6739__I1 mod.Data_Mem.F_M.MRAM\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5876_ _2099_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5247__S0 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7615_ _3747_ mod.Data_Mem.F_M.MRAM\[787\]\[1\] _3798_ _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4827_ mod.Data_Mem.F_M.src\[4\] _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8516__569 net569 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7247__I _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8595_ _0611_ net220 mod.Instr_Mem.instruction\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6364__A2 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6151__I _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4375__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5195__C _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7546_ _3731_ mod.Data_Mem.F_M.MRAM\[783\]\[7\] _3752_ _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4758_ _1421_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7477_ _3714_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4689_ _1226_ _1354_ _0997_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4127__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ _1937_ _1719_ _3035_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5875__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6359_ _2241_ _2244_ _2966_ _2969_ _1489_ _2784_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5627__A1 _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8029_ _0238_ net73 mod.Data_Mem.F_M.MRAM\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6978__I1 mod.Data_Mem.F_M.MRAM\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__A2 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4118__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__B _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5405__I _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5618__A1 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6437__S _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6830__A3 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout170_I net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout268_I net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3991_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5730_ _2158_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5661_ _2273_ _2123_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6346__A2 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7400_ _3673_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8002__CLK net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ _1197_ _1281_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8380_ _0476_ net120 mod.Data_Mem.F_M.MRAM\[784\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5592_ _1694_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7331_ _3603_ mod.Data_Mem.F_M.MRAM\[771\]\[0\] _3636_ _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4543_ _0635_ mod.Arithmetic.CN.I_in\[36\] _0893_ _0980_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4109__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7262_ _3593_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4474_ _1035_ _1036_ _1145_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _2105_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7193_ _3549_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _2757_ _2758_ _2759_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__A1 mod.Data_Mem.F_M.MRAM\[797\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5609__B2 mod.Data_Mem.F_M.MRAM\[796\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6075_ _1805_ _2690_ _2691_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5026_ _1541_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _3425_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ mod.Data_Mem.F_M.MRAM\[16\]\[4\] mod.Data_Mem.F_M.MRAM\[17\]\[4\] _2353_ _2549_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5859_ _2447_ _2481_ _1807_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6337__A2 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8578_ _0594_ net263 mod.Instr_Mem.instruction\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7529_ _3746_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5848__A1 _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5848__B2 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5225__I _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4520__A1 mod.Arithmetic.CN.I_in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6273__A1 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6025__A1 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8025__CLK net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__A2 _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8175__CLK net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7128__I1 mod.Data_Mem.F_M.MRAM\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5839__B2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6500__A2 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7551__S _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ _0825_ _0826_ _0675_ _0852_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_79_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4974__I _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout385_I net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__S _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7300__I1 mod.Data_Mem.F_M.MRAM\[768\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A2 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _3373_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7880_ _0106_ net170 mod.Data_Mem.F_M.MRAM\[26\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _3336_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4923__B _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ mod.Data_Mem.F_M.MRAM\[8\]\[4\] _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ _0645_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8501_ _0005_ net265 mod.Data_Mem.F_M.out_data\[77\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5713_ _2338_ mod.Data_Mem.F_M.MRAM\[28\]\[7\] _2311_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6693_ _3244_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6319__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8432_ _0528_ net192 mod.Data_Mem.F_M.MRAM\[792\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5644_ _2164_ _2275_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8363_ _0459_ net254 mod.Data_Mem.F_M.MRAM\[782\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4050__I0 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5575_ _2204_ _2205_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7314_ _3610_ _3626_ _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7819__A2 mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4526_ _1103_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8294_ _0390_ net91 mod.Data_Mem.F_M.MRAM\[772\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7245_ _3583_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4457_ _1127_ _1129_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4502__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _3543_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4388_ _0640_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__4884__I _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6127_ _2675_ _2741_ _2742_ _2080_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5058__A2 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__I0 mod.Data_Mem.F_M.MRAM\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _2674_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__I1 mod.Data_Mem.F_M.MRAM\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5009_ _1557_ _1636_ _1672_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6007__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4018__B1 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6558__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8198__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5369__I0 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5518__B1 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3963__I _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4995__S _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6494__A1 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5297__A2 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6495__B _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__I1 mod.Data_Mem.F_M.MRAM\[783\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7046__I0 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7349__I1 mod.Data_Mem.F_M.MRAM\[771\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7546__S _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout133_I net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4969__I _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6182__B1 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout300_I net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ mod.Data_Mem.F_M.MRAM\[5\]\[7\] mod.Data_Mem.F_M.MRAM\[4\]\[7\] _1878_ _2022_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4311_ _0898_ _0837_ _0897_ mod.Arithmetic.CN.I_in\[41\] _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5291_ mod.Data_Mem.F_M.MRAM\[769\]\[5\] _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__A1 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7030_ _3416_ mod.Data_Mem.F_M.MRAM\[18\]\[5\] _3457_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4242_ _0647_ mod.Arithmetic.ACTI.x\[2\] _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4173_ _0671_ _0846_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7080__I mod.Data_Mem.F_M.MRAM\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7285__I0 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7932_ _0158_ net377 mod.Data_Mem.F_M.MRAM\[8\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4799__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_490 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5460__A2 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7863_ _0089_ net382 mod.Data_Mem.F_M.MRAM\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8340__CLK net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ mod.Data_Mem.F_M.MRAM\[789\]\[2\] _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7908__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7794_ _3895_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6745_ _3273_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3957_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6676_ _3229_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8415_ _0511_ net88 mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8498__D _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5627_ _2259_ mod.Data_Mem.F_M.MRAM\[29\]\[0\] _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8346_ _0442_ net314 mod.Data_Mem.F_M.MRAM\[780\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ _2064_ mod.Data_Mem.F_M.MRAM\[30\]\[2\] mod.Data_Mem.F_M.MRAM\[31\]\[2\] _2196_
+ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ _1177_ _1179_ _1175_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8277_ _0373_ net111 mod.Data_Mem.F_M.MRAM\[770\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5489_ _1796_ mod.Data_Mem.F_M.MRAM\[31\]\[4\] _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__A1 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7228_ _3573_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7159_ _3248_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__I1 mod.Data_Mem.F_M.MRAM\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__I0 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3958__I _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5739__B1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6400__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5203__A2 _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4962__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4962__B2 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7165__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4190__A2 _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6467__A1 _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__A1 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__A2 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout250_I net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4860_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ mod.Arithmetic.CN.I_in\[23\] mod.Arithmetic.CN.I_in\[31\] _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6530_ _2261_ mod.Data_Mem.F_M.MRAM\[12\]\[6\] _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_119_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6461_ mod.Data_Mem.F_M.MRAM\[12\]\[2\] _1886_ _2525_ _2475_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8200_ _0085_ net11 net114 mod.I_addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__4705__A1 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5412_ _2070_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6392_ _2864_ _3001_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8131_ mod.Data_Mem.F_M.out_data\[41\] net52 net330 mod.Arithmetic.CN.I_in\[41\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_115_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5343_ mod.Data_Mem.F_M.MRAM\[791\]\[6\] mod.Data_Mem.F_M.MRAM\[788\]\[6\] mod.Data_Mem.F_M.MRAM\[789\]\[6\]
+ mod.Data_Mem.F_M.MRAM\[790\]\[6\] _1915_ _1917_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7803__I mod.Data_Mem.F_M.MRAM\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6458__A1 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8062_ _0271_ net80 mod.Data_Mem.F_M.MRAM\[20\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ mod.Data_Mem.F_M.MRAM\[788\]\[5\] _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ _3433_ _3446_ _3421_ _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4225_ _0897_ _0898_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5681__A2 mod.Data_Mem.F_M.MRAM\[29\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4156_ _0655_ _0824_ mod.Arithmetic.CN.I_in\[33\] _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_56_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4087_ _0734_ _0735_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7915_ _0141_ net368 mod.Data_Mem.F_M.MRAM\[10\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4383__B _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7846_ _3925_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3995__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7777_ _3885_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4989_ _1588_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _3267_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4944__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5926__C _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6659_ mod.Data_Mem.F_M.MRAM\[27\]\[1\] _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8236__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8329_ _0425_ net371 mod.Data_Mem.F_M.MRAM\[777\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7497__I0 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6449__A1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8386__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout340 net343 net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout351 net352 net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout362 net364 net362 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_120_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout373 net374 net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout384 net385 net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4880__B1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A1 _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6385__B1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5408__I _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4163__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5143__I _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4010_ mod.Arithmetic.I_out\[75\] _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_84_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5663__A2 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8109__CLK net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5961_ _2579_ mod.Data_Mem.F_M.MRAM\[5\]\[5\] _2580_ _2506_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7700_ mod.Data_Mem.F_M.MRAM\[793\]\[2\] _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4912_ _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3977__A2 mod.Arithmetic.CN.I_in\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5892_ _2510_ _2511_ _2512_ _2348_ _2513_ _2350_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_34_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7631_ _2043_ _3804_ _3809_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _1511_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7562_ _3767_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5974__I0 mod.Data_Mem.F_M.MRAM\[770\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _1435_ _1438_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_6513_ _2075_ mod.Data_Mem.F_M.MRAM\[0\]\[5\] _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7493_ _3711_ mod.Data_Mem.F_M.MRAM\[781\]\[3\] _3720_ _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6444_ _3051_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5351__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4154__A2 mod.Arithmetic.CN.I_in\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _2868_ _2037_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7533__I _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8114_ mod.Data_Mem.F_M.out_data\[24\] net46 net329 mod.Arithmetic.CN.I_in\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_115_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5326_ _1985_ _1986_ _1987_ _1988_ _1882_ _1666_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4378__B _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8045_ _0254_ net106 mod.Data_Mem.F_M.MRAM\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5257_ mod.Data_Mem.F_M.MRAM\[787\]\[4\] _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4208_ _0870_ _0872_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_111_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _1839_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4892__I _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ _0645_ _0811_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_29_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5957__A3 _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__A2 mod.Arithmetic.CN.I_in\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7829_ _3174_ _3909_ _3908_ _3915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4768__I1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6119__B1 _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4145__A2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3971__I _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5893__A2 _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout170 net171 net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_94_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout181 net183 net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout192 net194 net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_47_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4751__B _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5339__S _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7570__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4384__A2 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5581__B2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4042__I _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout213_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4490_ _1160_ _1082_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5074__S _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6160_ _1733_ _1715_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5111_ _1733_ _1777_ _1664_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6091_ _1501_ _1545_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6684__I1 mod.Data_Mem.F_M.MRAM\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5042_ _1517_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6993_ _3434_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6061__A2 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5944_ _2503_ mod.Data_Mem.F_M.MRAM\[14\]\[4\] _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5875_ _2056_ mod.Data_Mem.F_M.MRAM\[783\]\[3\] _2495_ _2496_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5247__S1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4826_ mod.Data_Mem.F_M.src\[2\] _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7614_ _3799_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8594_ _0610_ net115 mod.Instr_Mem.instruction\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7545_ _3756_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4375__A2 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4757_ _1422_ _1426_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7476_ _3615_ mod.Data_Mem.F_M.MRAM\[780\]\[4\] _3713_ _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4688_ _1353_ _1357_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6427_ _1767_ mod.Data_Mem.F_M.MRAM\[769\]\[1\] _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4887__I _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5875__A2 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6358_ mod.Data_Mem.F_M.MRAM\[781\]\[6\] _2745_ _2901_ mod.Data_Mem.F_M.MRAM\[780\]\[6\]
+ _2968_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_88_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _1966_ _1967_ _1970_ _1972_ _1698_ _1530_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6289_ _1525_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5627__A2 mod.Data_Mem.F_M.MRAM\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8028_ _0237_ net70 mod.Data_Mem.F_M.MRAM\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4571__B _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8574__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3966__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__C _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5563__A1 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5618__A2 mod.Data_Mem.F_M.MRAM\[797\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7615__I0 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6043__A2 mod.Data_Mem.F_M.MRAM\[19\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3990_ mod.Arithmetic.CN.F_in\[0\] _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout330_I net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6252__I _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ _2252_ mod.Data_Mem.F_M.MRAM\[28\]\[2\] _2254_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _1201_ _1258_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5591_ mod.Data_Mem.F_M.MRAM\[29\]\[4\] _2221_ _2222_ mod.Data_Mem.F_M.MRAM\[28\]\[4\]
+ _2227_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_128_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7330_ _3635_ _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4542_ _0636_ mod.Arithmetic.CN.I_in\[37\] _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7261_ mod.Data_Mem.F_M.MRAM\[31\]\[6\] _3319_ _3590_ _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5306__A1 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4473_ _1035_ _1036_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6212_ _2793_ _2799_ _2826_ _2367_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7192_ _3552_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _1740_ _1652_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout76_I net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6074_ mod.Data_Mem.F_M.MRAM\[13\]\[0\] _2083_ _2205_ mod.Data_Mem.F_M.MRAM\[12\]\[0\]
+ _2105_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_100_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5025_ _1692_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4293__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__A2 mod.Data_Mem.F_M.MRAM\[772\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _3393_ mod.Data_Mem.F_M.MRAM\[16\]\[1\] _3423_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__I0 _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5927_ _2395_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5793__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5858_ _2123_ _2444_ _2360_ _2479_ _2480_ _2168_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4809_ _1372_ _1380_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5545__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7194__S _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8577_ _0593_ net117 mod.Instr_Mem.instruction\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5789_ _2108_ _2412_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7528_ _3718_ mod.Data_Mem.F_M.MRAM\[783\]\[0\] _3745_ _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7459_ mod.Data_Mem.F_M.MRAM\[778\]\[6\] _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5950__B _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6025__A2 mod.Data_Mem.F_M.MRAM\[788\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6072__I _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4511__A2 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout280_I net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6247__I _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout378_I net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _3332_ _3298_ _3335_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6761_ _3287_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4578__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3973_ _0649_ mod.Arithmetic.CN.I_in\[24\] _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8500_ _0004_ net246 mod.Data_Mem.F_M.out_data\[76\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5712_ _2337_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6692_ _3243_ mod.Data_Mem.F_M.MRAM\[28\]\[2\] _3237_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8431_ _0527_ net90 mod.Data_Mem.F_M.MRAM\[791\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5643_ _2270_ _2272_ _2274_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8362_ _0458_ net292 mod.Data_Mem.F_M.MRAM\[782\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5574_ _2206_ _2176_ _2208_ _2211_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7313_ _3625_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4525_ _1159_ _1162_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8293_ _0389_ net143 mod.Data_Mem.F_M.MRAM\[772\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7244_ _3539_ mod.Data_Mem.F_M.MRAM\[30\]\[7\] _3579_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4456_ _1008_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4502__A2 mod.Arithmetic.CN.I_in\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7175_ mod.Data_Mem.F_M.MRAM\[22\]\[2\] _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4387_ _0956_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ _2182_ _2682_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__I1 mod.Data_Mem.F_M.MRAM\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6057_ _1693_ _2395_ _1535_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4266__A1 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7987__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _1675_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4018__A1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4018__B2 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6959_ _3413_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5945__B _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5518__A1 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5369__I1 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5518__B2 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6191__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5377__S0 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6494__A2 mod.Data_Mem.F_M.MRAM\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6067__I _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4257__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7046__I1 mod.Data_Mem.F_M.MRAM\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__C _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__A1 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8292__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 mod.Data_Mem.F_M.MRAM\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__B2 mod.Data_Mem.F_M.MRAM\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4310_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5290_ _1710_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4241_ _0648_ mod.Arithmetic.ACTI.x\[1\] _0669_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7361__I mod.Data_Mem.F_M.MRAM\[772\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__A1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4172_ _0669_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6237__A2 _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5296__I0 _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7931_ _0157_ net386 mod.Data_Mem.F_M.MRAM\[8\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5996__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4799__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_480 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_491 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7862_ _0088_ net378 mod.Data_Mem.F_M.MRAM\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5748__A1 _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6813_ _3325_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__I0 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout39_I net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7793_ _3312_ mod.Data_Mem.F_M.MRAM\[798\]\[4\] _3894_ _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _3278_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3956_ _0632_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4420__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ mod.Data_Mem.F_M.dest\[4\] mod.Data_Mem.F_M.dest\[2\] _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5626_ _2142_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8414_ _0510_ net87 mod.Data_Mem.F_M.MRAM\[788\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8345_ _0441_ net315 mod.Data_Mem.F_M.MRAM\[780\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5920__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5557_ _2094_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5056__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4508_ _1175_ _1177_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_8276_ _0372_ net110 mod.Data_Mem.F_M.MRAM\[770\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ _1840_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7227_ _3230_ _3464_ _3389_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4439_ _0644_ mod.Arithmetic.CN.I_in\[57\] _0922_ _1019_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7271__I mod.Data_Mem.F_M.MRAM\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7158_ _3532_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6109_ mod.Data_Mem.F_M.MRAM\[7\]\[0\] mod.Data_Mem.F_M.MRAM\[6\]\[0\] _2179_ _2726_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7089_ _3491_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4239__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8165__CLK net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5987__A1 _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__I1 mod.Data_Mem.F_M.MRAM\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5739__A1 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6787__I0 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5739__B2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4135__I _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__A2 mod.Data_Mem.F_M.MRAM\[780\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5675__B _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4962__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6164__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4190__A3 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6467__A2 mod.Data_Mem.F_M.MRAM\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8508__CLK net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6219__A2 _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4650__A1 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4045__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout243_I net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4790_ _1308_ _1315_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4402__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__S _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6260__I _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6460_ _3020_ _2479_ _3066_ _3063_ _1633_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5411_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6391_ _2866_ _2992_ _3000_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4705__A2 mod.Arithmetic.ACTI.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8130_ mod.Data_Mem.F_M.out_data\[40\] net51 net334 mod.Arithmetic.CN.I_in\[40\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5342_ _1872_ _2004_ _1863_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8061_ _0270_ net75 mod.Data_Mem.F_M.MRAM\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8136__RN net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ _1889_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7012_ _3388_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4224_ _0656_ _0835_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _0654_ _0830_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4086_ _0759_ _0761_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5969__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7914_ _0140_ net382 mod.Data_Mem.F_M.MRAM\[10\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4383__C _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7845_ mod.Data_Mem.F_M.MRAM\[9\]\[1\] _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7776_ _3806_ mod.Data_Mem.F_M.MRAM\[797\]\[5\] _3883_ _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4988_ _1641_ _1646_ _1654_ _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6727_ mod.Data_Mem.F_M.MRAM\[10\]\[6\] _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3939_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6658_ _3219_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7194__I0 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ mod.Data_Mem.F_M.MRAM\[797\]\[6\] _2221_ _1750_ mod.Data_Mem.F_M.MRAM\[796\]\[6\]
+ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6941__I0 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ _3184_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8328_ _0424_ net197 mod.Data_Mem.F_M.MRAM\[777\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8127__RN net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__A2 mod.Data_Mem.F_M.MRAM\[769\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7497__I1 mod.Data_Mem.F_M.MRAM\[781\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8259_ _0355_ net184 mod.Data_Mem.F_M.MRAM\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout330 net333 net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout341 net343 net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout352 net353 net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout363 net365 net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout374 net381 net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout385 net388 net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4880__A1 mod.Data_Mem.F_M.MRAM\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3969__I _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__C _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A1 mod.Data_Mem.F_M.MRAM\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__B2 mod.Data_Mem.F_M.MRAM\[12\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A3 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4699__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5424__I mod.Data_Mem.F_M.src\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout193_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__S _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__B1 mod.Data_Mem.F_M.MRAM\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout360_I net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6255__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5960_ _2464_ mod.Data_Mem.F_M.MRAM\[4\]\[5\] _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4911_ _1573_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5891_ mod.Data_Mem.F_M.MRAM\[2\]\[3\] mod.Data_Mem.F_M.MRAM\[3\]\[3\] _2420_ _2513_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7630_ _3322_ _3798_ _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6376__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ _1510_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7561_ _3725_ mod.Data_Mem.F_M.MRAM\[784\]\[4\] _3760_ _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4926__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4773_ _1440_ _1439_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7086__I mod.Data_Mem.F_M.MRAM\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5974__I1 mod.Data_Mem.F_M.MRAM\[771\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6512_ _2689_ mod.Data_Mem.F_M.MRAM\[12\]\[5\] _3115_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7492_ _3723_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _3040_ _3050_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6374_ _2713_ _2982_ _2983_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7628__A1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5325_ mod.Data_Mem.F_M.MRAM\[3\]\[6\] mod.Data_Mem.F_M.MRAM\[2\]\[6\] _1890_ _1988_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8113_ mod.Data_Mem.F_M.out_data\[23\] net40 net274 mod.Arithmetic.CN.I_in\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__7750__S _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4378__C _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8044_ _0253_ net78 mod.Data_Mem.F_M.MRAM\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5256_ _1694_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _0880_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4311__B1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ _1845_ mod.Data_Mem.F_M.MRAM\[771\]\[3\] _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4138_ _0650_ _0813_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4069_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4614__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5002__C _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7828_ _3914_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7759_ _3782_ mod.Data_Mem.F_M.MRAM\[796\]\[6\] _3872_ _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6119__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4393__A3 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6119__B2 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6914__I0 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout160 net161 net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_94_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout171 net174 net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout182 net183 net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout193 net194 net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__A1 mod.Data_Mem.F_M.MRAM\[781\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6358__B2 mod.Data_Mem.F_M.MRAM\[780\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5419__I _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6905__I0 _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6530__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _1774_ mod.Data_Mem.F_M.MRAM\[769\]\[2\] _1776_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _1648_ _1605_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _1705_ _1707_ _1708_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4439__A4 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _3433_ _3371_ _3421_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5943_ _2562_ mod.Data_Mem.F_M.MRAM\[5\]\[4\] _2563_ _2510_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5874_ _2202_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout21_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _3771_ mod.Data_Mem.F_M.MRAM\[787\]\[0\] _3798_ _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4825_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8376__CLK net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8593_ _0609_ net226 mod.Instr_Mem.instruction\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7544_ _3729_ mod.Data_Mem.F_M.MRAM\[783\]\[6\] _3752_ _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4756_ mod.Arithmetic.CN.I_in\[39\] _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7475_ _3706_ _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4687_ _1353_ _1356_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6426_ _2309_ mod.Data_Mem.F_M.MRAM\[781\]\[1\] _2374_ _3033_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6521__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6357_ _2746_ _2967_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5064__I _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ mod.Data_Mem.F_M.MRAM\[3\]\[5\] mod.Data_Mem.F_M.MRAM\[2\]\[5\] _1971_ _1972_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _1546_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5999__I _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8027_ _0236_ net70 mod.Data_Mem.F_M.MRAM\[16\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _1514_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_76_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4571__C _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3982__I _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6512__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7893__CLK net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8249__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7615__I1 mod.Data_Mem.F_M.MRAM\[787\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout156_I net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7565__S _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6200__B1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4053__I mod.Arithmetic.CN.I_in\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout323_I net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _1201_ _1258_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5590_ _2223_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4541_ _1209_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7260_ _3592_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6503__A1 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4472_ _1039_ _1144_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5306__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7551__I0 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6211_ _2219_ _2814_ _2819_ _2825_ _2737_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_7191_ _3527_ mod.Data_Mem.F_M.MRAM\[29\]\[1\] _3550_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _1602_ _1650_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7303__I0 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6708__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6073_ _2689_ mod.Data_Mem.F_M.MRAM\[14\]\[0\] mod.Data_Mem.F_M.MRAM\[15\]\[0\] _2506_
+ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4817__A1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _1522_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout69_I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__B1 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6975_ _3424_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7782__A3 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5926_ _2359_ _2546_ _2098_ _2440_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_81_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5793__A2 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5857_ mod.Data_Mem.F_M.MRAM\[16\]\[2\] mod.Data_Mem.F_M.MRAM\[17\]\[2\] _2337_ _2480_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5059__I _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4808_ _0625_ _1367_ _1368_ _1381_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_8576_ _0592_ net263 mod.Instr_Mem.instruction\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7790__I0 _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5788_ _2410_ _1686_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4898__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ _3744_ _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4739_ _1335_ _1343_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7458_ _3702_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6111__C _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7542__I0 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6409_ _3016_ mod.Data_Mem.F_M.MRAM\[13\]\[0\] _2375_ _3017_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7389_ mod.Data_Mem.F_M.MRAM\[774\]\[3\] _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5950__C _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5856__I0 mod.Data_Mem.F_M.MRAM\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4808__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__A1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8541__CLK net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6281__I0 mod.Data_Mem.F_M.MRAM\[789\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4587__A3 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__A1 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8071__CLK net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4511__A3 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5432__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5472__A1 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout273_I net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6760_ mod.Data_Mem.F_M.MRAM\[8\]\[3\] _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6972__A1 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5711_ _1639_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6691_ _3242_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8430_ _0526_ net91 mod.Data_Mem.F_M.MRAM\[791\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5642_ _2273_ _2121_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8361_ _0457_ net293 mod.Data_Mem.F_M.MRAM\[782\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6212__B _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5573_ _2209_ mod.Data_Mem.F_M.MRAM\[30\]\[3\] _2210_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7312_ _3622_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4524_ _1165_ _1187_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__7524__I0 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8292_ _0388_ net95 mod.Data_Mem.F_M.MRAM\[772\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7243_ _3582_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4455_ _0614_ mod.Arithmetic.ACTI.x\[4\] _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4386_ _0640_ mod.Arithmetic.CN.I_in\[20\] _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7174_ _3542_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4502__A3 mod.Arithmetic.CN.I_in\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ _2165_ _2739_ _2740_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _2523_ _2656_ _2673_ _2407_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5007_ _1674_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _3397_ mod.Data_Mem.F_M.MRAM\[15\]\[3\] _3409_ _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5909_ mod.Data_Mem.F_M.MRAM\[784\]\[4\] mod.Data_Mem.F_M.MRAM\[785\]\[4\] _2516_
+ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6889_ mod.Data_Mem.F_M.MRAM\[4\]\[4\] _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7507__A3 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5518__A2 mod.Data_Mem.F_M.MRAM\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5369__I2 _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8559_ _0063_ net275 mod.Data_Mem.F_M.out_data\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6122__B _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__I _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8094__CLK net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7515__I0 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5377__S1 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__I _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7931__CLK net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5454__A1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4257__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5206__A1 _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5509__A2 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6182__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__I _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4193__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout119_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__I1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4240_ _0641_ mod.Arithmetic.CN.I_in\[66\] _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__A1 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4496__A2 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout390_I net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4171_ _0668_ mod.Arithmetic.ACTI.x\[1\] _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5296__I1 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7930_ _0156_ net171 mod.Data_Mem.F_M.MRAM\[8\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_470 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5996__A2 mod.Data_Mem.F_M.MRAM\[772\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_481 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_492 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_7861_ _3917_ _3919_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__A1 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__B _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6812_ mod.Data_Mem.F_M.MRAM\[789\]\[1\] _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7792_ _3888_ _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__I1 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _3246_ mod.Data_Mem.F_M.MRAM\[0\]\[3\] _3274_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4956__B1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3955_ _0614_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4420__A2 mod.Arithmetic.CN.I_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6674_ _3227_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8413_ _0509_ net139 mod.Data_Mem.F_M.MRAM\[788\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5625_ _2069_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6173__A2 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8344_ _0440_ net312 mod.Data_Mem.F_M.MRAM\[780\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5556_ _2194_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5920__A2 mod.Data_Mem.F_M.MRAM\[773\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6369__S _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4507_ _0646_ _1178_ _1064_ _1070_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8275_ _0371_ net183 mod.Data_Mem.F_M.MRAM\[770\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5487_ _2112_ _2127_ _2130_ _2132_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7954__CLK net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7226_ _3572_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4438_ _1109_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5684__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__I _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7157_ _3531_ mod.Data_Mem.F_M.MRAM\[12\]\[3\] _3525_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4369_ _0952_ _0975_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ mod.Data_Mem.F_M.MRAM\[1\]\[0\] _1539_ _1813_ mod.Data_Mem.F_M.MRAM\[0\]\[0\]
+ _2702_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7088_ mod.Data_Mem.F_M.MRAM\[21\]\[7\] _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ mod.Data_Mem.F_M.MRAM\[16\]\[7\] mod.Data_Mem.F_M.MRAM\[17\]\[7\] _2420_ _2657_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5987__A2 mod.Data_Mem.F_M.MRAM\[786\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6832__S _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__C1 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5739__A2 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8090__RN net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4175__A1 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5911__A2 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3990__I mod.Arithmetic.CN.F_in\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5675__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6806__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5817__I3 mod.Data_Mem.F_M.MRAM\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3989__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5358__S _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4402__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout236_I net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4061__I _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _2059_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4166__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6390_ _2865_ _2999_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4996__I _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5341_ _2000_ _2001_ _2002_ _2003_ _1911_ _1591_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_86_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__S _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8060_ _0269_ net89 mod.Data_Mem.F_M.MRAM\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5272_ _1698_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4469__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7011_ _3227_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4223_ mod.Arithmetic.CN.I_in\[42\] _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4154_ _0635_ mod.Arithmetic.CN.I_in\[33\] _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4085_ _0760_ _0714_ _0727_ _0728_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5620__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5969__A2 mod.Data_Mem.F_M.MRAM\[782\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6091__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7913_ _0139_ net155 mod.Data_Mem.F_M.MRAM\[10\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_fanout51_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4641__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7748__S _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7844_ _3924_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7775_ _3884_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _1559_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6726_ _3266_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3938_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6657_ mod.Data_Mem.F_M.MRAM\[27\]\[0\] _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6146__A2 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7194__I1 mod.Data_Mem.F_M.MRAM\[29\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ _1708_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6588_ mod.I_addr\[6\] _3183_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8327_ _0423_ net192 mod.Data_Mem.F_M.MRAM\[776\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5539_ _1695_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7282__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8258_ _0354_ net149 mod.Data_Mem.F_M.MRAM\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7209_ _3523_ mod.Data_Mem.F_M.MRAM\[2\]\[0\] _3562_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout320 net322 net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_8189_ _0299_ net196 mod.Data_Mem.F_M.MRAM\[19\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout331 net332 net331 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout342 net343 net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout353 net367 net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout364 net365 net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout375 net376 net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout386 net388 net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__4880__A2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8282__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6082__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6385__A2 _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__B1 mod.Data_Mem.F_M.MRAM\[798\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6932__I1 mod.Data_Mem.F_M.MRAM\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4699__A2 mod.Arithmetic.CN.I_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6696__I0 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6737__S _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout186_I net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5440__I _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__B2 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4084__B1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout353_I net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4910_ _1566_ _1572_ _1578_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ mod.Data_Mem.F_M.MRAM\[18\]\[3\] mod.Data_Mem.F_M.MRAM\[19\]\[3\] _2427_ _2512_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4841_ _1503_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6376__A2 _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4387__A1 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8005__CLK net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7560_ _3766_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4772_ mod.Arithmetic.CN.I_in\[55\] _1441_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6204__C _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6511_ _2374_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7491_ _3640_ mod.Data_Mem.F_M.MRAM\[781\]\[2\] _3720_ _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4139__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6442_ _3044_ _3046_ _3048_ _3049_ _2080_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5887__A1 _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__CLK net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _2889_ _2035_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8112_ mod.Data_Mem.F_M.out_data\[22\] net40 net274 mod.Arithmetic.CN.I_in\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7628__A2 _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5324_ mod.Data_Mem.F_M.MRAM\[1\]\[6\] mod.Data_Mem.F_M.MRAM\[0\]\[6\] _1878_ _1987_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout99_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8043_ _0252_ net71 mod.Data_Mem.F_M.MRAM\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ _1732_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6300__A2 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4206_ _0878_ _0874_ _0876_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_87_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4311__B2 mod.Arithmetic.CN.I_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5186_ _1604_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4137_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _0680_ _0683_ _0700_ _0706_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_56_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5811__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4614__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7827_ _3908_ _3913_ _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7277__I mod.Data_Mem.F_M.MRAM\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4378__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7758_ _3874_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6114__C _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6709_ _3256_ mod.Data_Mem.F_M.MRAM\[28\]\[6\] _3250_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7316__A1 _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6119__A2 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7689_ _3838_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4393__A4 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6914__I1 mod.Data_Mem.F_M.MRAM\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5461__S _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4302__A1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout150 net151 net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout161 net165 net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout172 net173 net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout183 net215 net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout194 net199 net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6055__A1 _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8028__CLK net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7555__A1 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__A2 _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6305__B _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4369__A1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6905__I1 mod.Data_Mem.F_M.MRAM\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6530__A2 mod.Data_Mem.F_M.MRAM\[12\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout101_I net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4541__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6294__B2 mod.Data_Mem.F_M.MRAM\[12\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5341__I0 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _1574_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__B _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6266__I _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6046__A1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6991_ _3234_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7298__S _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6841__I0 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5942_ _2503_ mod.Data_Mem.F_M.MRAM\[4\]\[4\] _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_94_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5873_ _2261_ mod.Data_Mem.F_M.MRAM\[782\]\[3\] _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_90_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7612_ _3797_ _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4824_ _1492_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8592_ _0608_ net220 mod.Instr_Mem.instruction\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7543_ _3755_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout14_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4755_ mod.Arithmetic.CN.I_in\[37\] _1423_ _1214_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4080__I0 mod.Arithmetic.CN.I_in\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4780__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6506__C1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7474_ _3712_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4686_ _0618_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_49_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6425_ _2353_ mod.Data_Mem.F_M.MRAM\[780\]\[1\] _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6521__A2 mod.Data_Mem.F_M.MRAM\[780\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6356_ _2268_ mod.Data_Mem.F_M.MRAM\[783\]\[6\] mod.Data_Mem.F_M.MRAM\[782\]\[6\]
+ _2904_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ _1511_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6287_ _1537_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5281__S _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8026_ _0235_ net209 mod.Data_Mem.F_M.MRAM\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5332__I0 mod.Data_Mem.F_M.MRAM\[17\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6285__B2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _1902_ _1702_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _1511_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5080__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6037__A1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__I0 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5260__A2 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8470__CLK net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4771__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6512__A2 mod.Data_Mem.F_M.MRAM\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4287__B1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5204__B _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6028__A1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6814__I mod.Data_Mem.F_M.MRAM\[789\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6750__S _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout149_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__A1 _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6200__B2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5366__S _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout316_I net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4540_ _1210_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7000__I0 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4471_ _1042_ _1046_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6503__A2 mod.Data_Mem.F_M.MRAM\[769\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6210_ _1899_ _2824_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4514__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7190_ _3551_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _2700_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7303__I1 mod.Data_Mem.F_M.MRAM\[768\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5314__I0 mod.Data_Mem.F_M.MRAM\[19\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _2271_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5023_ _1681_ mod.Data_Mem.F_M.MRAM\[789\]\[1\] _1690_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6019__B2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5490__A2 mod.Data_Mem.F_M.MRAM\[30\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6974_ _3386_ mod.Data_Mem.F_M.MRAM\[16\]\[0\] _3423_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5925_ mod.Data_Mem.F_M.MRAM\[18\]\[4\] mod.Data_Mem.F_M.MRAM\[19\]\[4\] _2353_ _2546_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8493__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5856_ mod.Data_Mem.F_M.MRAM\[14\]\[2\] mod.Data_Mem.F_M.MRAM\[15\]\[2\] _1774_ _2479_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4807_ _1325_ _1475_ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8575_ _0079_ net245 mod.Data_Mem.F_M.out_data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5787_ _2304_ mod.Data_Mem.F_M.MRAM\[787\]\[1\] _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7790__I1 mod.Data_Mem.F_M.MRAM\[798\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7526_ _3407_ _3705_ _3387_ _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4738_ _1208_ _1210_ _1338_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7457_ mod.Data_Mem.F_M.MRAM\[778\]\[5\] _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4669_ mod.Arithmetic.CN.I_in\[46\] _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7542__I1 mod.Data_Mem.F_M.MRAM\[783\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7491__S _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4505__A1 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _2500_ mod.Data_Mem.F_M.MRAM\[12\]\[0\] _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7388_ _3667_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ _2883_ _2946_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5803__I _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6258__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8009_ _0218_ net305 mod.Data_Mem.F_M.MRAM\[14\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5856__I1 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5481__A2 _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__B1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5233__A2 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6430__A1 _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4992__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7465__I _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6733__A2 mod.Data_Mem.F_M.dest\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8501__D _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4744__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6497__A1 _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4347__I1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6249__A1 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5472__A2 mod.Data_Mem.F_M.MRAM\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout266_I net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7576__S _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5710_ _2309_ mod.Data_Mem.F_M.MRAM\[29\]\[7\] _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6690_ net5 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7221__I0 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5641_ _1916_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7375__I mod.Data_Mem.F_M.MRAM\[773\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8360_ _0456_ net287 mod.Data_Mem.F_M.MRAM\[782\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4735__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ _2063_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6212__C _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7311_ _3624_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8291_ _0387_ net139 mod.Data_Mem.F_M.MRAM\[772\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5824__S _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7524__I1 mod.Data_Mem.F_M.MRAM\[782\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6488__A1 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7242_ _3537_ mod.Data_Mem.F_M.MRAM\[30\]\[6\] _3579_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _0642_ mod.Arithmetic.ACTI.x\[3\] _0915_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7173_ mod.Data_Mem.F_M.MRAM\[22\]\[1\] _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4385_ _0616_ _0697_ mod.Arithmetic.CN.I_in\[19\] _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout81_I net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6124_ mod.Data_Mem.F_M.MRAM\[781\]\[1\] _2193_ _2195_ mod.Data_Mem.F_M.MRAM\[780\]\[1\]
+ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_112_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _2520_ _2665_ _2672_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5006_ _1673_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _3412_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7883__CLK net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5908_ _2395_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6888_ _3366_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5839_ _2431_ _2124_ _2459_ _2396_ _2461_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6176__B1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8239__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__B2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8558_ _0062_ net275 mod.Data_Mem.F_M.out_data\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7509_ _3718_ mod.Data_Mem.F_M.MRAM\[782\]\[0\] _3734_ _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8489_ _0585_ net140 mod.Data_Mem.F_M.MRAM\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6479__A1 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5961__C _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5454__A2 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3988__I mod.Arithmetic.ACTI.x\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5206__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6403__A1 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6403__B2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5201__C _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4265__I0 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5909__S _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__I0 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8231__D mod.P1.instr_reg\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5693__A2 mod.Data_Mem.F_M.MRAM\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4170_ _0668_ mod.Arithmetic.CN.I_in\[65\] _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout383_I net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5296__I2 _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_460 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_471 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_482 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6274__I _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7860_ _3917_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xtiny_user_project_493 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_51_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _3324_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7791_ _3893_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5819__S _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _3277_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4956__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ _0623_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__B2 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6673_ net3 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8412_ _0508_ net85 mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5624_ _2092_ _2256_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8343_ _0439_ net156 mod.Data_Mem.F_M.MRAM\[778\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8531__CLK net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5555_ _1546_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4506_ mod.Arithmetic.CN.I_in\[29\] _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8274_ _0370_ net203 mod.Data_Mem.F_M.MRAM\[770\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5486_ _2066_ _2131_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7225_ _3539_ mod.Data_Mem.F_M.MRAM\[2\]\[7\] _3567_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4437_ _0993_ _0999_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5684__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7156_ _3245_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4368_ _0902_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_63_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _2722_ mod.Data_Mem.F_M.MRAM\[3\]\[0\] _1808_ _2723_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7087_ _3490_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4299_ _0722_ _0820_ _0884_ _0715_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_58_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5436__A2 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6038_ _2409_ _2648_ _2655_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6117__C _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6397__B1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5729__S _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7989_ mod.Instr_Mem.instruction\[22\] net11 net100 mod.Data_Mem.F_M.src\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6397__C2 _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6492__S0 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6149__B1 mod.Data_Mem.F_M.MRAM\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5528__I _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5372__A1 mod.Data_Mem.F_M.MRAM\[783\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3989__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6822__I mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout131_I net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout229_I net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4166__A2 mod.Arithmetic.CN.I_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__S _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5340_ mod.Data_Mem.F_M.MRAM\[775\]\[6\] mod.Data_Mem.F_M.MRAM\[774\]\[6\] _1831_
+ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5271_ mod.Data_Mem.F_M.MRAM\[799\]\[5\] _1934_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7010_ _3444_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4222_ _0634_ mod.Arithmetic.CN.I_in\[42\] _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4153_ _0828_ mod.Arithmetic.CN.I_in\[48\] _0674_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4084_ _0756_ _0757_ _0714_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_95_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4517__I mod.Arithmetic.CN.I_in\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6091__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7912_ _0138_ net205 mod.Data_Mem.F_M.MRAM\[10\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout44_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7843_ mod.Data_Mem.F_M.MRAM\[9\]\[0\] _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6732__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5977__I0 mod.Data_Mem.F_M.MRAM\[786\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7774_ _3778_ mod.Data_Mem.F_M.MRAM\[797\]\[4\] _3883_ _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4986_ _1648_ _1650_ _1653_ _1617_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6725_ mod.Data_Mem.F_M.MRAM\[10\]\[5\] _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3937_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5729__I0 mod.Data_Mem.F_M.MRAM\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6656_ _3218_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _2229_ mod.Data_Mem.F_M.MRAM\[799\]\[6\] mod.Data_Mem.F_M.MRAM\[798\]\[6\]
+ _1816_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4157__A2 _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _3178_ mod.I_addr\[5\] _3179_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5354__B2 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8326_ _0422_ net382 mod.Data_Mem.F_M.MRAM\[776\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _1575_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5106__A1 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8257_ _0353_ net149 mod.Data_Mem.F_M.MRAM\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5083__I _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5469_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7208_ _3561_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5657__A2 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8188_ _0298_ net195 mod.Data_Mem.F_M.MRAM\[19\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout310 net325 net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout321 net322 net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout332 net333 net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout343 net352 net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7139_ _3508_ mod.Data_Mem.F_M.MRAM\[19\]\[5\] _3518_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout354 net356 net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout365 net366 net365 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout376 net380 net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout387 net388 net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_100_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5032__B _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8577__CLK net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4396__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__B2 _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5258__I _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6217__S0 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6310__C _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6696__I1 mod.Data_Mem.F_M.MRAM\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4320__A2 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5721__I _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A2 mod.Data_Mem.F_M.MRAM\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout179_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7648__I mod.Data_Mem.F_M.MRAM\[790\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout346_I net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7944__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4387__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _1354_ mod.Arithmetic.CN.I_in\[54\] _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7584__S _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6510_ _2579_ mod.Data_Mem.F_M.MRAM\[13\]\[5\] _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7490_ _3722_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5336__A1 mod.Data_Mem.F_M.MRAM\[783\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6441_ _2105_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6372_ _2887_ _2036_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6220__C _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8111_ mod.Data_Mem.F_M.out_data\[21\] net43 net278 mod.Arithmetic.CN.I_in\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5323_ mod.Data_Mem.F_M.MRAM\[7\]\[6\] mod.Data_Mem.F_M.MRAM\[6\]\[6\] _1876_ _1986_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8042_ _0251_ net195 mod.Data_Mem.F_M.MRAM\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5254_ _1703_ _1918_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4205_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4311__A2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5631__I _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ mod.Data_Mem.F_M.MRAM\[770\]\[3\] _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4136_ _0615_ mod.Arithmetic.CN.I_in\[25\] _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A2 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4247__I mod.Arithmetic.CN.I_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7558__I _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7826_ mod.I_addr\[3\] _3911_ _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__A1 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7757_ _3806_ mod.Data_Mem.F_M.MRAM\[796\]\[5\] _3872_ _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4969_ _1567_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6708_ _3255_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7688_ mod.Data_Mem.F_M.MRAM\[792\]\[4\] _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7316__A2 _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ mod.Data_Mem.F_M.MRAM\[26\]\[7\] _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8309_ _0405_ net158 mod.Data_Mem.F_M.MRAM\[774\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout140 net141 net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout151 net152 net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout162 net165 net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout173 net174 net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout184 net186 net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout195 net196 net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7967__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7555__A2 _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6515__B1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6748__S _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout296_I net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5341__I1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5451__I _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4495__C _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7618__I0 _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__A2 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4057__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6990_ _3432_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6841__I1 mod.Data_Mem.F_M.MRAM\[769\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5941_ _2207_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5099__S _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6282__I _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5872_ _2415_ _2130_ _2486_ _2493_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7611_ _3296_ _3604_ _3758_ _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4823_ mod.Data_Mem.F_M.src\[1\] _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8122__CLK net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8591_ _0607_ net385 mod.Data_Mem.F_M.MRAM\[9\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7542_ _3754_ mod.Data_Mem.F_M.MRAM\[783\]\[5\] _3752_ _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4754_ _1185_ _1423_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4080__I1 mod.Arithmetic.I_out\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7473_ _3711_ mod.Data_Mem.F_M.MRAM\[780\]\[3\] _3707_ _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6506__B1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6231__B _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4685_ mod.Arithmetic.CN.I_in\[54\] _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5626__I _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6506__C2 _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4530__I mod.Arithmetic.CN.I_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8272__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6424_ _3019_ _2430_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6109__I0 mod.Data_Mem.F_M.MRAM\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6355_ mod.Data_Mem.F_M.MRAM\[13\]\[6\] _2900_ _2194_ mod.Data_Mem.F_M.MRAM\[12\]\[6\]
+ _2965_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_89_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5306_ _1711_ _1968_ _1969_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _2876_ _2882_ _2892_ _2898_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6285__A2 _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8025_ _0234_ net301 mod.Data_Mem.F_M.MRAM\[16\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5237_ mod.Data_Mem.F_M.MRAM\[783\]\[4\] _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5332__I1 mod.Data_Mem.F_M.MRAM\[16\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4296__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__I0 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _1830_ _1832_ _1833_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7489__S _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4119_ _0792_ _0791_ _0795_ mod.Arithmetic.ACTI.x\[6\] _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _1764_ _1765_ _1568_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6832__I1 mod.Data_Mem.F_M.MRAM\[769\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7288__I _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5310__B _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7809_ mod.Data_Mem.F_M.MRAM\[7\]\[4\] _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5548__A1 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6920__I _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5536__I _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4287__A1 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6028__A2 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5787__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8145__CLK net361 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5220__B _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__A2 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4211__A1 mod.Arithmetic.CN.I_in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout211_I net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7000__I1 mod.Data_Mem.F_M.MRAM\[17\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout309_I net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4470_ _1047_ _1084_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4514__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6140_ _2177_ _2754_ _2755_ _2710_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7464__A1 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ _2677_ _2681_ _1728_ _2687_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5314__I1 mod.Data_Mem.F_M.MRAM\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__B1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5022_ _1570_ _1689_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6019__A2 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6973_ _3422_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6941__S _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ _2409_ _2534_ _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5855_ _2346_ _2477_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _1328_ _1386_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8574_ _0078_ net264 mod.Data_Mem.F_M.out_data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4202__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5786_ _2179_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7525_ _3743_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5950__A1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4737_ _1350_ _1362_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5356__I _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7456_ _3701_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4668_ _1203_ mod.Arithmetic.CN.I_in\[45\] _0984_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6407_ _2590_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4505__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6750__I0 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5702__A1 _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7387_ mod.Data_Mem.F_M.MRAM\[774\]\[2\] _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7571__I _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4599_ _1261_ _1262_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6338_ _2771_ _2947_ _2948_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6258__A2 _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6269_ _2877_ _2879_ _2880_ _2881_ _2072_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5091__I _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8008_ _0217_ net302 mod.Data_Mem.F_M.MRAM\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A3 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8168__CLK net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__C1 _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A1 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__B2 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7998__RN net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4441__A1 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4744__A2 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__I _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8175__RN net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6741__I0 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4680__A1 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6046__B _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout161_I net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7989__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3970_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout259_I net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5480__I0 mod.Data_Mem.F_M.MRAM\[30\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6185__A1 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _2271_ mod.Data_Mem.F_M.MRAM\[796\]\[1\] _2262_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5232__I0 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5571_ _2054_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6980__I0 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5932__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4735__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7310_ _3603_ mod.Data_Mem.F_M.MRAM\[770\]\[0\] _3623_ _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4522_ _1188_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_129_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _0386_ net185 mod.Data_Mem.F_M.MRAM\[772\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8166__RN net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7241_ _3581_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4453_ mod.Arithmetic.CN.I_in\[65\] _1012_ _0643_ mod.Arithmetic.ACTI.x\[2\] _1126_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5904__I _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7172_ _3541_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4384_ _1054_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ _2611_ mod.Data_Mem.F_M.MRAM\[783\]\[1\] mod.Data_Mem.F_M.MRAM\[782\]\[1\]
+ _2085_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _2557_ _2667_ _2669_ _2671_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ mod.Data_Mem.F_M.src\[8\] _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4671__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7767__S _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4255__I mod.Arithmetic.CN.I_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6956_ _3395_ mod.Data_Mem.F_M.MRAM\[15\]\[2\] _3409_ _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5907_ _2056_ mod.Data_Mem.F_M.MRAM\[788\]\[4\] _2527_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6887_ mod.Data_Mem.F_M.MRAM\[4\]\[3\] _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6176__A1 mod.Data_Mem.F_M.MRAM\[781\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5838_ _2418_ _1788_ _2419_ _2460_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6176__B2 mod.Data_Mem.F_M.MRAM\[780\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6403__C _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4726__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5923__A1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8557_ _0061_ net280 mod.Data_Mem.F_M.out_data\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5769_ _2387_ _2097_ _2390_ _2393_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7508_ _3733_ _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8488_ _0584_ net164 mod.Data_Mem.F_M.MRAM\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6479__A2 mod.Data_Mem.F_M.MRAM\[769\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8157__RN net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7439_ mod.Data_Mem.F_M.MRAM\[777\]\[4\] _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7007__S _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__A1 _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6100__B2 _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4662__A1 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__A1 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6403__A2 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4414__A1 _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5611__B1 mod.Data_Mem.F_M.MRAM\[30\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7203__I1 mod.Data_Mem.F_M.MRAM\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5214__I0 mod.Data_Mem.F_M.MRAM\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5925__S _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8333__CLK net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8148__RN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout376_I net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5599__C _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5296__I3 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_450 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_461 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_472 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_483 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_494 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__S _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6810_ mod.Data_Mem.F_M.MRAM\[789\]\[0\] _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4405__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7790_ _3309_ mod.Data_Mem.F_M.MRAM\[798\]\[3\] _3889_ _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__B1 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6741_ _3243_ mod.Data_Mem.F_M.MRAM\[0\]\[2\] _3274_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3953_ mod.Arithmetic.CN.I_in\[8\] _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4956__A2 mod.Data_Mem.F_M.MRAM\[799\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6504__B _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__I _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6672_ _3226_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8411_ _0507_ net142 mod.Data_Mem.F_M.MRAM\[788\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5623_ _2085_ _2097_ _2251_ _2255_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_8342_ _0438_ net385 mod.Data_Mem.F_M.MRAM\[778\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5554_ _1538_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4505_ _0958_ _1176_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8273_ _0369_ net203 mod.Data_Mem.F_M.MRAM\[770\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6705__I0 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5485_ _1761_ _2069_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7224_ _3571_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4436_ _0930_ _0995_ _0996_ _0997_ _0994_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_63_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7155_ _3530_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4367_ _0970_ _0974_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6106_ _2571_ mod.Data_Mem.F_M.MRAM\[2\]\[0\] _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7086_ mod.Data_Mem.F_M.MRAM\[21\]\[6\] _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7130__I0 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5436__A3 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6037_ _2535_ _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7497__S _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A1 _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7988_ mod.Instr_Mem.instruction\[17\] net21 net226 mod.P1.instr_reg\[17\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6397__B2 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6939_ _3399_ mod.Data_Mem.F_M.MRAM\[14\]\[4\] _3400_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6492__S1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_161_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6149__A1 _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6944__I0 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6321__A1 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6321__B2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5480__S _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4635__A1 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3989__A3 mod.Arithmetic.CN.I_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6388__A1 mod.Data_Mem.F_M.MRAM\[781\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6388__B2 mod.Data_Mem.F_M.MRAM\[780\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5719__I _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6935__I0 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout124_I net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6560__A1 _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _1597_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6312__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5115__A2 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4221_ _0893_ _0894_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4152_ _0817_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7112__I0 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4083_ _0713_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7911_ _0137_ net368 mod.Data_Mem.F_M.MRAM\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7842_ _3923_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7110__S _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout37_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7773_ _3877_ _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5977__I1 mod.Data_Mem.F_M.MRAM\[787\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__I _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _1588_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6724_ _3265_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3936_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6926__I0 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5729__I1 mod.Data_Mem.F_M.MRAM\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6655_ mod.Data_Mem.F_M.MRAM\[25\]\[7\] _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5606_ mod.Data_Mem.F_M.MRAM\[29\]\[6\] _2082_ _2222_ mod.Data_Mem.F_M.MRAM\[28\]\[6\]
+ _2240_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6551__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _3182_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8325_ _0421_ net166 mod.Data_Mem.F_M.MRAM\[776\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ _1642_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8256_ _0352_ net163 mod.Data_Mem.F_M.MRAM\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6303__A1 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5106__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5468_ _2115_ _1627_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7207_ _3270_ _3272_ _3389_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout300 net310 net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4419_ _0894_ _0980_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8187_ _0297_ net196 mod.Data_Mem.F_M.MRAM\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout311 net312 net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5399_ _1673_ _2059_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout322 net324 net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout333 net338 net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7138_ _3519_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout344 net347 net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout355 net360 net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout366 net367 net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6409__B _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout377 net378 net377 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout388 net389 net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _3481_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5539__I _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5593__A2 mod.Data_Mem.F_M.MRAM\[799\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4396__A3 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6217__S1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7754__I _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6542__A1 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7590__I0 _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7896__CLK net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7342__I0 _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4320__A3 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__I mod.Arithmetic.CN.I_in\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4084__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5449__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5033__A1 mod.Data_Mem.F_M.MRAM\[799\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout241_I net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout339_I net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _0624_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__I mod.Data_Mem.F_M.MRAM\[791\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6440_ _3047_ _2282_ _3008_ _2443_ _2450_ _2484_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5336__A2 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6533__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6371_ _2893_ _2979_ _2980_ _2897_ _2072_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8110_ mod.Data_Mem.F_M.out_data\[20\] net42 net278 mod.Arithmetic.CN.I_in\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5322_ mod.Data_Mem.F_M.MRAM\[5\]\[6\] mod.Data_Mem.F_M.MRAM\[4\]\[6\] _1874_ _1985_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6297__B1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8041_ _0250_ net195 mod.Data_Mem.F_M.MRAM\[18\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5253_ mod.Data_Mem.F_M.MRAM\[791\]\[4\] mod.Data_Mem.F_M.MRAM\[788\]\[4\] mod.Data_Mem.F_M.MRAM\[789\]\[4\]
+ mod.Data_Mem.F_M.MRAM\[790\]\[4\] _1915_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__8051__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4956__C _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5895__I0 mod.Data_Mem.F_M.MRAM\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4204_ _0874_ _0876_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5184_ _1591_ _1843_ _1849_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6229__B _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8525__564 net564 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4135_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6944__S _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ mod.Arithmetic.CN.I_in\[14\] _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7013__A2 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7825_ _3907_ _3912_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__B1 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7756_ _3873_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__A2 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4968_ _1633_ _1634_ _1635_ mod.Data_Mem.F_M.MRAM\[15\]\[1\] _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6707_ net9 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7687_ _3837_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5295__S _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4899_ _1567_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6638_ _3209_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5327__A2 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6524__A1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7572__I0 _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6569_ _0612_ _3169_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5094__I _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8308_ _0404_ net79 mod.Data_Mem.F_M.MRAM\[774\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7324__I0 _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8239_ _0335_ net132 mod.Data_Mem.F_M.MRAM\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7015__S _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4838__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout130 net131 net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout141 net146 net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout152 net153 net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout163 net164 net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout174 net175 net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout185 net186 net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout196 net198 net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6055__A3 _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__B _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5263__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5269__I _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7484__I _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4901__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6515__A1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7563__I0 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__B2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6321__C _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8074__CLK net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout191_I net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4057__A2 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__A1 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5940_ _2558_ mod.Data_Mem.F_M.MRAM\[2\]\[4\] _2559_ _2560_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _2488_ _2489_ _2491_ _2492_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4083__I _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7610_ _3796_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4822_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8590_ _0606_ net193 mod.Data_Mem.F_M.MRAM\[9\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7541_ _3315_ _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4753_ mod.Arithmetic.CN.I_in\[38\] _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6512__B _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6004__S _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6506__A1 _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7472_ _3308_ _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6506__B2 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4684_ mod.Arithmetic.CN.I_in\[52\] _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ _3030_ _2275_ _3023_ _2412_ _2417_ _3022_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__6939__S _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7306__I0 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6354_ _2902_ _2964_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8567__CLK net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _1906_ mod.Data_Mem.F_M.MRAM\[0\]\[5\] _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6285_ _2893_ _2894_ _2896_ _2897_ _1899_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8024_ _0233_ net301 mod.Data_Mem.F_M.MRAM\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5236_ _1871_ _1885_ _1887_ _1898_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7609__I1 mod.Data_Mem.F_M.MRAM\[786\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _1529_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5798__B _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4118_ _0744_ _0784_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ mod.Data_Mem.F_M.MRAM\[773\]\[2\] mod.Data_Mem.F_M.MRAM\[772\]\[2\] _1763_
+ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7569__I _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ _0716_ _0718_ _0725_ _0630_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7808_ _3902_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7793__I0 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7739_ _3863_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4220__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8097__CLK net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5484__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4287__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5787__A2 mod.Data_Mem.F_M.MRAM\[787\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5928__S _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7784__I0 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4211__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7536__I0 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6051__C _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout204_I net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5462__I _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6070_ _2083_ _2683_ _2686_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A1 _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ mod.Data_Mem.F_M.MRAM\[788\]\[1\] _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5475__B2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6972_ _3269_ _3270_ _3421_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6226__C _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5923_ _2535_ _2543_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5854_ _2440_ _2474_ _2475_ _2360_ _2476_ _2444_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_61_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4805_ _1328_ _1386_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8573_ _0077_ net282 mod.Data_Mem.F_M.out_data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5785_ _2371_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4202__A2 mod.Arithmetic.CN.I_in\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7524_ _3731_ mod.Data_Mem.F_M.MRAM\[782\]\[7\] _3739_ _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4736_ _1294_ _1402_ _1405_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5950__A2 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3961__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7455_ mod.Data_Mem.F_M.MRAM\[778\]\[4\] _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4667_ _1252_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7957__CLK net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6406_ _2861_ _3007_ _3014_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7386_ _3666_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5702__A2 mod.Data_Mem.F_M.MRAM\[29\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6750__I1 mod.Data_Mem.F_M.MRAM\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4598_ mod.Arithmetic.ACTI.x\[6\] _1268_ _0802_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6337_ _1582_ _2000_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6268_ _2833_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8007_ _0216_ net301 mod.Data_Mem.F_M.MRAM\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4917__S _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5219_ _1560_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6199_ _2806_ _2813_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6415__B1 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6415__C2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6430__A3 _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6281__I3 mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__I0 mod.Data_Mem.F_M.MRAM\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4441__A2 mod.Arithmetic.CN.I_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6931__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7518__I0 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6741__I1 mod.Data_Mem.F_M.MRAM\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6329__S0 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8112__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7203__S _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4680__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7002__I _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8262__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6501__S0 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4968__B1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5480__I1 mod.Data_Mem.F_M.MRAM\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout154_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7757__I0 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6185__A2 mod.Data_Mem.F_M.MRAM\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5457__I _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout321_I net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7509__I0 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _2207_ mod.Data_Mem.F_M.MRAM\[31\]\[3\] _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6980__I1 mod.Data_Mem.F_M.MRAM\[16\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4521_ _1190_ _1079_ _1191_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4991__I0 mod.Data_Mem.F_M.MRAM\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7240_ _3569_ mod.Data_Mem.F_M.MRAM\[30\]\[5\] _3579_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5145__B1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4452_ _0667_ mod.Arithmetic.CN.I_in\[68\] _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5696__A1 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6288__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7171_ mod.Data_Mem.F_M.MRAM\[22\]\[0\] _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4383_ _0643_ _0959_ _0813_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6122_ _2688_ _2697_ _2738_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5448__A1 _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _2555_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5004_ _1656_ _1670_ _1671_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_fanout67_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6237__B _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__I mod.Arithmetic.CN.I_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4671__A2 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6952__S _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _3411_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4423__A2 mod.Arithmetic.CN.I_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5906_ _2526_ mod.Data_Mem.F_M.MRAM\[789\]\[4\] _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6886_ _3365_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7748__I0 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ _2420_ mod.Data_Mem.F_M.MRAM\[789\]\[2\] _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6176__A2 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8556_ _0060_ net277 mod.Data_Mem.F_M.out_data\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5923__A2 _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5768_ _2391_ mod.Data_Mem.F_M.MRAM\[788\]\[0\] _2392_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7507_ _3634_ _3387_ _3389_ _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4982__I0 mod.Data_Mem.F_M.MRAM\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _1274_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8487_ _0583_ net102 mod.Data_Mem.F_M.MRAM\[798\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5699_ _2277_ _2140_ _2324_ _2326_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7438_ _3692_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5687__A1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7369_ mod.Data_Mem.F_M.MRAM\[773\]\[1\] _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8285__CLK net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__A2 _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8093__RN net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5611__A1 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5611__B2 _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A2 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5214__I1 mod.Data_Mem.F_M.MRAM\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6836__I _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_440 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__B _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_451 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4653__A2 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5850__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_462 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_473 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_fanout369_I net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_484 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_495 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__A1 mod.Data_Mem.F_M.MRAM\[797\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6571__I mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5602__B2 mod.Data_Mem.F_M.MRAM\[796\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ _3276_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3952_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output8_I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6671_ mod.Data_Mem.F_M.MRAM\[27\]\[7\] _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8410_ _0506_ net190 mod.Data_Mem.F_M.MRAM\[788\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4169__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5622_ _2252_ mod.Data_Mem.F_M.MRAM\[796\]\[0\] _2254_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8341_ _0437_ net371 mod.Data_Mem.F_M.MRAM\[778\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5553_ mod.Data_Mem.F_M.MRAM\[797\]\[2\] _2176_ _2189_ mod.Data_Mem.F_M.MRAM\[796\]\[2\]
+ _2191_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7108__S _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4504_ _0613_ _1062_ mod.Arithmetic.CN.I_in\[29\] _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8272_ _0368_ net187 mod.Data_Mem.F_M.MRAM\[770\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5484_ _2128_ mod.Data_Mem.F_M.MRAM\[799\]\[3\] _2129_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6705__I1 mod.Data_Mem.F_M.MRAM\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5669__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7223_ _3537_ mod.Data_Mem.F_M.MRAM\[2\]\[6\] _3567_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5136__B _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6947__S _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4435_ _1000_ _1001_ _1106_ _1107_ _1004_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_132_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7154_ _3529_ mod.Data_Mem.F_M.MRAM\[12\]\[2\] _3525_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4366_ _0951_ _1037_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6105_ _1783_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7085_ _3489_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7130__I1 mod.Data_Mem.F_M.MRAM\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4297_ _0618_ mod.Arithmetic.CN.I_in\[11\] _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__A1 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _2415_ _2649_ _2650_ _2454_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_100_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7987_ mod.Instr_Mem.instruction\[13\] net16 net219 mod.P1.instr_reg\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6397__A2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8075__RN net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6938_ _3390_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ mod.Data_Mem.F_M.MRAM\[6\]\[2\] _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6944__I1 mod.Data_Mem.F_M.MRAM\[14\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8539_ _0043_ net277 mod.Data_Mem.F_M.out_data\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7018__S _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6321__A2 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4332__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4635__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5832__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8523__D _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8300__CLK net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6935__I1 mod.Data_Mem.F_M.MRAM\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__A1 _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5735__I _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4571__A1 mod.Arithmetic.CN.I_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout117_I net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6312__A2 _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4220_ _0824_ _0830_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4323__A1 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5520__B1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ _0825_ _0826_ _0675_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7112__I1 mod.Data_Mem.F_M.MRAM\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4082_ _0756_ _0757_ _0710_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_95_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7910_ _0136_ net308 mod.Data_Mem.F_M.MRAM\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7841_ _0610_ _3922_ _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7772_ _3882_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4984_ mod.Data_Mem.F_M.MRAM\[1\]\[1\] mod.Data_Mem.F_M.MRAM\[0\]\[1\] _1651_ _1652_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6723_ mod.Data_Mem.F_M.MRAM\[10\]\[4\] _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3935_ mod.Arithmetic.CN.F_in\[0\] _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _3217_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6926__I1 mod.Data_Mem.F_M.MRAM\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _2223_ _2239_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6585_ mod.I_addr\[5\] _3181_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6551__A2 mod.Data_Mem.F_M.MRAM\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5645__I _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8324_ _0420_ net205 mod.Data_Mem.F_M.MRAM\[776\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5536_ _2082_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8255_ _0351_ net116 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _2114_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6303__A2 _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7206_ _3560_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5362__I0 _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5511__B1 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4418_ _0619_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8186_ _0296_ net191 mod.Data_Mem.F_M.MRAM\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout301 net304 net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _2058_ _1534_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xfanout312 net319 net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout323 net324 net323 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7137_ _3456_ mod.Data_Mem.F_M.MRAM\[19\]\[4\] _3518_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout334 net336 net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _0992_ _1002_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_101_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout345 net347 net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout356 net360 net356 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout367 net390 net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout378 net380 net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout389 net390 net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7068_ mod.Data_Mem.F_M.MRAM\[20\]\[5\] _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5814__A1 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _2635_ _2636_ _2637_ _2555_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7319__A1 _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4396__A4 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6542__A2 mod.Data_Mem.F_M.MRAM\[768\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5555__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7342__I1 mod.Data_Mem.F_M.MRAM\[771\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5290__I _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5805__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7211__S _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6230__A1 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5033__A2 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout234_I net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4792__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7030__I0 _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6533__A2 mod.Data_Mem.F_M.MRAM\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__A1 mod.Arithmetic.CN.I_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _2029_ _2030_ _2895_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5321_ mod.Data_Mem.F_M.MRAM\[15\]\[6\] _1679_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6297__A1 mod.Data_Mem.F_M.MRAM\[781\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8040_ _0249_ net195 mod.Data_Mem.F_M.MRAM\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6297__B2 mod.Data_Mem.F_M.MRAM\[780\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5252_ _1916_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5895__I1 mod.Data_Mem.F_M.MRAM\[15\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4203_ _0809_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5183_ _1844_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6049__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8346__CLK net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4065_ _0738_ _0736_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7549__A1 _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8163__D mod.Data_Mem.F_M.out_data\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7824_ _3907_ _3911_ _3912_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8496__CLK net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6221__A1 _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__B2 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7755_ _3778_ mod.Data_Mem.F_M.MRAM\[796\]\[4\] _3872_ _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4967_ _1619_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5575__A3 _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6706_ _3254_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7686_ mod.Data_Mem.F_M.MRAM\[792\]\[3\] _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5980__B1 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4898_ _1524_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7021__I0 _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6637_ mod.Data_Mem.F_M.MRAM\[26\]\[6\] _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6524__A2 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6568_ mod.I_addr\[1\] _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8307_ _0403_ net161 mod.Data_Mem.F_M.MRAM\[774\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5519_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7324__I1 mod.Data_Mem.F_M.MRAM\[770\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6499_ _1623_ _3103_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8238_ _0334_ net107 mod.Data_Mem.F_M.MRAM\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4838__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout120 net130 net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_8169_ mod.Data_Mem.F_M.out_data\[79\] net27 net264 mod.Arithmetic.I_out\[79\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout131 net136 net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout142 net144 net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout153 net154 net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout164 net165 net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout175 net176 net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout186 net189 net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout197 net198 net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6934__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6460__B2 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8073__D mod.P3.Res\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7563__I1 mod.Data_Mem.F_M.MRAM\[784\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__A1 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5341__I3 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout184_I net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5254__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout351_I net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _2369_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6203__A1 _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _1489_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7540_ _3753_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4752_ _0622_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7003__I0 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7471_ _3710_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4683_ mod.Arithmetic.CN.I_in\[53\] _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6506__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _2090_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6353_ _2903_ mod.Data_Mem.F_M.MRAM\[15\]\[6\] mod.Data_Mem.F_M.MRAM\[14\]\[6\] _2253_
+ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5190__A1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7306__I1 mod.Data_Mem.F_M.MRAM\[768\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5304_ mod.Data_Mem.F_M.MRAM\[1\]\[5\] _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6284_ _2833_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8023_ _0232_ net210 mod.Data_Mem.F_M.MRAM\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5235_ _1899_ _1629_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5493__A2 mod.Data_Mem.F_M.MRAM\[798\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ mod.Data_Mem.F_M.MRAM\[791\]\[3\] mod.Data_Mem.F_M.MRAM\[790\]\[3\] _1831_
+ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4117_ _0747_ _0772_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5097_ mod.Data_Mem.F_M.MRAM\[775\]\[2\] mod.Data_Mem.F_M.MRAM\[774\]\[2\] _1763_
+ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6442__B2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4048_ _0691_ _0724_ _0708_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7886__CLK net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7786__S _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7242__I0 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7807_ mod.Data_Mem.F_M.MRAM\[7\]\[3\] _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5999_ _2617_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7793__I1 mod.Data_Mem.F_M.MRAM\[798\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4756__A1 mod.Arithmetic.CN.I_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7738_ mod.Data_Mem.F_M.MRAM\[795\]\[5\] _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7669_ _3828_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5181__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5054__B _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5484__A2 mod.Data_Mem.F_M.MRAM\[799\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6808__I0 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6433__A1 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__C _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7233__I0 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7784__I1 mod.Data_Mem.F_M.MRAM\[798\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8531__D _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4211__A3 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7536__I1 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6121__B1 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A2 _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5020_ _1681_ mod.Data_Mem.F_M.MRAM\[787\]\[1\] _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5899__B _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6424__A1 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6971_ _3420_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5922_ _2415_ _2536_ _2537_ _2454_ _2542_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4986__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ mod.Data_Mem.F_M.MRAM\[18\]\[2\] mod.Data_Mem.F_M.MRAM\[19\]\[2\] _1796_ _2476_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6523__B _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4738__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4822__I _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4804_ _1406_ _1432_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8572_ _0076_ net247 mod.Data_Mem.F_M.out_data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5784_ _2408_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout12_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7523_ _3742_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _0625_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8534__CLK net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7454_ _3700_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3961__A2 mod.Arithmetic.CN.I_in\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4666_ mod.Arithmetic.CN.I_in\[46\] _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4978__B _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _2108_ _2380_ _3012_ _3013_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5163__A1 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7385_ mod.Data_Mem.F_M.MRAM\[774\]\[1\] _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4597_ mod.P2.Rout_reg\[0\] _0678_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6336_ _1569_ _2001_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6267_ _1895_ _1894_ _1896_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8006_ _0215_ net233 mod.Data_Mem.F_M.MRAM\[13\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5218_ _1875_ _1877_ _1879_ _1881_ _1882_ _1666_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_57_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6198_ _2674_ _2809_ _2812_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7207__A3 _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5149_ _1504_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6415__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__B2 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7215__I0 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6018__I1 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6152__C _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7518__I1 mod.Data_Mem.F_M.MRAM\[782\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6329__S1 _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6406__A1 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__S1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__B2 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8557__CLK net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7757__I1 mod.Data_Mem.F_M.MRAM\[796\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4196__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7509__I1 mod.Data_Mem.F_M.MRAM\[782\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout314_I net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4520_ mod.Arithmetic.CN.I_in\[11\] _1078_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4991__I1 mod.Data_Mem.F_M.MRAM\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ _1008_ _1014_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5145__A1 mod.Data_Mem.F_M.MRAM\[22\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5696__A2 mod.Data_Mem.F_M.MRAM\[797\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7170_ _3540_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4382_ _0668_ mod.Arithmetic.CN.I_in\[26\] _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ _1728_ _2721_ _2729_ _2736_ _2737_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__A2 mod.Data_Mem.F_M.MRAM\[798\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ mod.Data_Mem.F_M.MRAM\[14\]\[7\] mod.Data_Mem.F_M.MRAM\[15\]\[7\] _2320_ _2670_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _1555_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _3393_ mod.Data_Mem.F_M.MRAM\[15\]\[1\] _3409_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5905_ _2400_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__I _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6885_ mod.Data_Mem.F_M.MRAM\[4\]\[2\] _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5836_ _2296_ _1797_ _2458_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7924__CLK net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8555_ _0059_ net328 mod.Data_Mem.F_M.out_data\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5767_ _1774_ mod.Data_Mem.F_M.MRAM\[789\]\[0\] _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7506_ _3732_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4718_ _1277_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4982__I1 mod.Data_Mem.F_M.MRAM\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8486_ _0582_ net102 mod.Data_Mem.F_M.MRAM\[798\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5698_ _2325_ mod.Data_Mem.F_M.MRAM\[796\]\[5\] _2084_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7437_ mod.Data_Mem.F_M.MRAM\[777\]\[3\] _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4649_ _1307_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4501__B _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5687__A2 mod.Data_Mem.F_M.MRAM\[796\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _3657_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6319_ _2772_ _1940_ _2930_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7299_ _3616_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5611__A2 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4178__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7773__I _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A1 _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4637__I _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_430 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_441 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_452 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_463 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_474 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_485 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_496 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7052__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout264_I net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5989__I0 mod.Data_Mem.F_M.MRAM\[784\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__A2 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3951_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6670_ _3225_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5621_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4169__A2 _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6563__B1 _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8340_ _0436_ net205 mod.Data_Mem.F_M.MRAM\[778\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5552_ _1648_ _2190_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4503_ _1173_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5118__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8271_ _0367_ net127 mod.Data_Mem.F_M.MRAM\[768\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5483_ _1792_ mod.Data_Mem.F_M.MRAM\[798\]\[3\] _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5669__A2 mod.Data_Mem.F_M.MRAM\[28\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7222_ _3570_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4434_ _1016_ _1021_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7153_ _3242_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4365_ _0948_ _1025_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7124__S _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6104_ _2183_ _2712_ _2720_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7084_ mod.Data_Mem.F_M.MRAM\[21\]\[5\] _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _0965_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7291__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6035_ _2538_ _2651_ _2652_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7986_ mod.Instr_Mem.instruction\[11\] net16 net219 mod.P1.instr_reg\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6937_ _3248_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6868_ _3356_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8102__CLK net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5357__A1 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ mod.Data_Mem.F_M.MRAM\[18\]\[1\] mod.Data_Mem.F_M.MRAM\[19\]\[1\] _2337_ _2443_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7593__I _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6799_ _3315_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8538_ _0042_ net346 mod.Data_Mem.F_M.out_data\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5327__B _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5109__A1 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8469_ _0565_ net235 mod.Data_Mem.F_M.MRAM\[796\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8252__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5841__I _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5596__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5596__B2 _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__S _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5899__A2 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6113__S _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5952__S _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5520__A1 mod.Data_Mem.F_M.MRAM\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4323__A2 mod.Arithmetic.CN.I_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5751__I _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4150_ _0654_ _0657_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout381_I net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6783__S _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4081_ _0630_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6320__I0 _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7678__I mod.Data_Mem.F_M.MRAM\[791\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7840_ _0080_ _3171_ _3921_ _3916_ _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7771_ _3309_ mod.Data_Mem.F_M.MRAM\[797\]\[3\] _3878_ _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4983_ _1542_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6722_ _3264_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3934_ _0612_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6653_ mod.Data_Mem.F_M.MRAM\[25\]\[6\] _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6531__B _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4830__I _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ _1747_ mod.Data_Mem.F_M.MRAM\[31\]\[6\] mod.Data_Mem.F_M.MRAM\[30\]\[6\] _2166_
+ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8275__CLK net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6584_ _3178_ _3179_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8323_ _0419_ net370 mod.Data_Mem.F_M.MRAM\[776\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6958__S _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5535_ _2154_ _2131_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8254_ _0350_ net116 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5466_ _1916_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7205_ _3539_ mod.Data_Mem.F_M.MRAM\[29\]\[7\] _3549_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4417_ mod.Arithmetic.CN.I_in\[36\] _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5511__A1 _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8185_ _0295_ net107 mod.Data_Mem.F_M.MRAM\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5362__I1 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5511__B2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5397_ _1502_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout302 net304 net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_67_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout313 net319 net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_67_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout324 net325 net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7136_ _3512_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4348_ _1004_ _1016_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_86_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout335 net336 net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout346 net347 net346 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout357 net359 net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout368 net369 net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_7067_ _3480_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout379 net380 net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4279_ _0693_ _0810_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ mod.Data_Mem.F_M.MRAM\[14\]\[6\] mod.Data_Mem.F_M.MRAM\[15\]\[6\] _2582_ _2637_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5578__A1 _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7969_ _0195_ net163 mod.Data_Mem.F_M.MRAM\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4250__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7319__A2 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5057__B _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5772__S _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5502__A1 _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__C1 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8148__CLK net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4851__S _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6230__A2 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8298__CLK net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4241__A1 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__I0 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5746__I _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7030__I1 mod.Data_Mem.F_M.MRAM\[18\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout227_I net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5041__I0 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4544__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5741__A1 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5320_ _1900_ _1964_ _1983_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6297__A2 _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _1504_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4202_ _0641_ mod.Arithmetic.CN.I_in\[18\] _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5182_ _1845_ mod.Data_Mem.F_M.MRAM\[773\]\[3\] _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4097__I mod.Arithmetic.ACTI.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6049__A2 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4133_ _0632_ mod.Arithmetic.CN.I_in\[17\] _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4064_ _0729_ _0734_ _0735_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_68_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__I _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6018__S _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7823_ _3171_ _3908_ _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__S _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6221__A2 mod.Data_Mem.F_M.MRAM\[14\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7754_ _3866_ _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4966_ mod.Data_Mem.F_M.MRAM\[31\]\[1\] _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4232__A1 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6705_ _3253_ mod.Data_Mem.F_M.MRAM\[28\]\[5\] _3250_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7685_ _3836_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6261__B _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__A1 _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__B2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6636_ _3208_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6688__S _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _3083_ _3158_ _3160_ _3168_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_69_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8306_ _0402_ net190 mod.Data_Mem.F_M.MRAM\[774\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5518_ _2157_ mod.Data_Mem.F_M.MRAM\[30\]\[0\] mod.Data_Mem.F_M.MRAM\[31\]\[0\] _2158_
+ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6498_ _3058_ _2549_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8237_ _0333_ net132 mod.Data_Mem.F_M.MRAM\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5391__I _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ _1535_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4299__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4299__B2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout110 net112 net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout121 net124 net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_8168_ mod.Data_Mem.F_M.out_data\[78\] net27 net266 mod.Arithmetic.I_out\[78\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_2
XFILLER_59_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout132 net134 net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout143 net144 net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7119_ _3252_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout154 net178 net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__4936__S _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout165 net176 net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout176 net177 net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_8099_ mod.Data_Mem.F_M.out_data\[9\] net52 net344 mod.Arithmetic.CN.I_in\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5099__I0 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout187 net189 net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_74_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6445__C1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout198 net199 net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_47_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5343__S0 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5799__A1 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5799__B2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A2 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5971__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4774__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5566__I _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5326__I1 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__B1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6346__B _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout177_I net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4462__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4820_ mod.Data_Mem.F_M.src\[8\] _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout344_I net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A1 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4751_ _1203_ mod.Arithmetic.CN.I_in\[46\] _1209_ _1340_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7470_ _3640_ mod.Data_Mem.F_M.MRAM\[780\]\[2\] _3707_ _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4682_ mod.Arithmetic.CN.I_in\[61\] _1135_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8196__RN net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6421_ _3015_ _3029_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5714__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6352_ _2950_ _2953_ _2959_ _2962_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8313__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ mod.Data_Mem.F_M.MRAM\[7\]\[5\] mod.Data_Mem.F_M.MRAM\[6\]\[5\] _1682_ _1967_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6283_ _1925_ _1926_ _2895_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5478__B1 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8022_ _0231_ net122 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _1674_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5165_ _1768_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4116_ _0787_ _0786_ _0791_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5096_ _1710_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4047_ mod.Arithmetic.I_out\[72\] _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6442__A2 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6770__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7242__I1 mod.Data_Mem.F_M.MRAM\[30\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7806_ _3901_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5998_ _1757_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7737_ _3862_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5953__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _1614_ _1616_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7668_ mod.Data_Mem.F_M.MRAM\[791\]\[2\] _3828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6619_ mod.Data_Mem.F_M.MRAM\[24\]\[5\] _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5705__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7599_ _3612_ _3789_ _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4893__C _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6418__C1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6808__I1 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5316__S0 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7630__A1 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A2 mod.Data_Mem.F_M.MRAM\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7233__I1 mod.Data_Mem.F_M.MRAM\[30\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__I0 mod.Data_Mem.F_M.MRAM\[769\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5944__A1 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5899__C _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout294_I net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8102__RN net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6791__S _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6970_ mod.Data_Mem.F_M.dest\[4\] _3372_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5921_ _2538_ _2539_ _2541_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4986__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ mod.Data_Mem.F_M.MRAM\[2\]\[2\] mod.Data_Mem.F_M.MRAM\[3\]\[2\] _1786_ _2475_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ _1444_ _1452_ _1472_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5935__A1 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4738__A2 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8571_ _0075_ net334 mod.Data_Mem.F_M.out_data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6983__I0 _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _2073_ _2365_ _2367_ _2405_ _2407_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_7522_ _3729_ mod.Data_Mem.F_M.MRAM\[782\]\[6\] _3739_ _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4734_ mod.Arithmetic.CN.I_in\[63\] _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7453_ mod.Data_Mem.F_M.MRAM\[778\]\[3\] _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3961__A3 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4665_ _1202_ mod.Arithmetic.CN.I_in\[45\] _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5934__I _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6031__S _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6404_ _2098_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7384_ _3665_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5163__A2 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ _0805_ _0859_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6966__S _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6335_ _2842_ _2944_ _2945_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6112__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6266_ _2878_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _0214_ net259 mod.Data_Mem.F_M.MRAM\[13\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5217_ _1647_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4674__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6197_ _1643_ _2810_ _2811_ _2767_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5871__B1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5602__C _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ mod.Data_Mem.F_M.MRAM\[6\]\[3\] _1608_ _1812_ _1813_ _1560_ _1814_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__S _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4285__I _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8209__CLK net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5079_ _1607_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4426__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7596__I _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7215__I1 mod.Data_Mem.F_M.MRAM\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8359__CLK net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6974__I0 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6351__A1 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__B2 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8079__D mod.P3.Res\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7151__I0 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6103__A1 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4665__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5614__B1 mod.Data_Mem.F_M.MRAM\[798\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4968__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4798__C _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout307_I net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6342__A1 _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4450_ _1009_ _1013_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5145__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6342__B2 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7876__CLK net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4381_ _0957_ _0960_ _0961_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_98_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ _2359_ _2189_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _2562_ mod.Data_Mem.F_M.MRAM\[5\]\[7\] _2668_ _2510_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _1660_ _1665_ _1667_ _1669_ _1619_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4408__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _3410_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8501__CLK net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5929__I _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4833__I _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5904_ _2432_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6026__S _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6884_ _3364_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5835_ _2325_ mod.Data_Mem.F_M.MRAM\[785\]\[2\] _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6030__B1 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8554_ _0058_ net342 mod.Data_Mem.F_M.out_data\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6581__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _1840_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7505_ _3731_ mod.Data_Mem.F_M.MRAM\[781\]\[7\] _3726_ _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4717_ _1280_ _1283_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8485_ _0581_ net110 mod.Data_Mem.F_M.MRAM\[798\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5697_ _1747_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ _3691_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6333__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4648_ _1174_ _1310_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6696__S _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7367_ mod.Data_Mem.F_M.MRAM\[773\]\[0\] _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4579_ mod.Arithmetic.CN.I_in\[61\] _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4895__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6318_ _1737_ _1941_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7298_ _3615_ mod.Data_Mem.F_M.MRAM\[768\]\[4\] _3606_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6249_ _2861_ _2862_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8031__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4647__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7320__S _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6947__I0 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A2 _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4886__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7124__I0 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7824__A1 _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8537__D _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4638__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_420 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_121_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_431 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_442 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_453 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_464 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_475 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_486 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_497 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7052__A2 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3950_ mod.P2.Rout_reg\[0\] mod.P2.Rout_reg\[1\] _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout257_I net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5620_ _1493_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6563__A1 mod.Data_Mem.F_M.MRAM\[780\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _1954_ mod.Data_Mem.F_M.MRAM\[799\]\[2\] mod.Data_Mem.F_M.MRAM\[798\]\[2\]
+ _2088_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4502_ _0639_ mod.Arithmetic.CN.I_in\[21\] mod.Arithmetic.CN.I_in\[20\] _1174_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8270_ _0366_ net127 mod.Data_Mem.F_M.MRAM\[768\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6315__A1 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _2094_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7221_ _3569_ mod.Data_Mem.F_M.MRAM\[2\]\[5\] _3567_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4433_ _1004_ _1016_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8054__CLK net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7152_ _3528_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4364_ _0976_ _1024_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6103_ _2685_ _2716_ _2719_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7083_ _3488_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4295_ _0966_ _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A1 _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7291__A2 _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout72_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _2378_ mod.Data_Mem.F_M.MRAM\[772\]\[7\] _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7985_ mod.Instr_Mem.instruction\[10\] net18 net218 mod.P1.instr_reg\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5054__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _3398_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4801__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6929__I0 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6867_ mod.Data_Mem.F_M.MRAM\[6\]\[1\] _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ mod.Data_Mem.F_M.MRAM\[2\]\[1\] mod.Data_Mem.F_M.MRAM\[3\]\[1\] _1786_ _2442_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5357__A2 _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6554__A1 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6798_ net8 _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8537_ _0041_ net344 mod.Data_Mem.F_M.out_data\[33\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5749_ _2373_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8468_ _0564_ net236 mod.Data_Mem.F_M.MRAM\[796\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7419_ mod.Data_Mem.F_M.MRAM\[776\]\[2\] _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8399_ _0495_ net104 mod.Data_Mem.F_M.MRAM\[786\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4096__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__A1 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7050__S _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A1 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5348__A2 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6545__B2 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8077__CLK net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7345__I0 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7225__S _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4859__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5520__A2 _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4080_ mod.Arithmetic.CN.I_in\[17\] mod.Arithmetic.I_out\[73\] _0709_ _0757_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6320__I1 _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5284__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout374_I net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7770_ _3881_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4982_ mod.Data_Mem.F_M.MRAM\[3\]\[1\] mod.Data_Mem.F_M.MRAM\[2\]\[1\] _1649_ _1650_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6721_ mod.Data_Mem.F_M.MRAM\[10\]\[3\] _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3933_ mod.I_addr\[0\] _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _3216_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7584__I0 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__A1 _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5603_ _2220_ _2235_ _2238_ _2218_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6583_ _3180_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8322_ _0418_ net370 mod.Data_Mem.F_M.MRAM\[776\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5534_ _2174_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8253_ _0349_ net116 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5465_ _2093_ _2097_ _2103_ _2113_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4986__C _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7204_ _3559_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4416_ _0982_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8184_ _0294_ net76 mod.Data_Mem.F_M.MRAM\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5511__A2 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5396_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout303 net304 net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5163__B _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6974__S _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7135_ _3517_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout314 net318 net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_114_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout325 net326 net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4347_ _1018_ _1019_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout336 net337 net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout347 net351 net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout358 net359 net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout369 net374 net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7066_ mod.Data_Mem.F_M.MRAM\[20\]\[4\] _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4278_ _0883_ _0886_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5275__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6472__B1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ mod.Data_Mem.F_M.MRAM\[2\]\[6\] mod.Data_Mem.F_M.MRAM\[3\]\[6\] _2075_ _2636_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7968_ _0194_ net140 mod.Data_Mem.F_M.MRAM\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _3385_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7899_ _0125_ net197 mod.Data_Mem.F_M.MRAM\[27\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_168_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6527__A1 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6013__I _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5889__I0 mod.Data_Mem.F_M.MRAM\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5502__A2 mod.Data_Mem.F_M.MRAM\[31\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6463__B1 _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__C2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4241__A2 mod.Arithmetic.ACTI.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__I _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__A1 _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__I1 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__C _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5248__B _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5963__S _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5041__I1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout122_I net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5741__A2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ _1543_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_64_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ mod.Arithmetic.CN.I_in\[24\] _0813_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5181_ _1604_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4132_ _0631_ _0652_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4063_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A1 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7822_ mod.I_addr\[0\] _3169_ _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout35_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7753_ _3871_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4965_ _1622_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5937__I _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6704_ _3252_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__A1 _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7684_ mod.Data_Mem.F_M.MRAM\[792\]\[2\] _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5980__A2 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4896_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6635_ mod.Data_Mem.F_M.MRAM\[26\]\[5\] _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _2861_ _3162_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4997__B _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8305_ _0401_ net170 mod.Data_Mem.F_M.MRAM\[774\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5517_ _2114_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6497_ _3096_ _3097_ _3101_ _2106_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5672__I _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8236_ _0332_ net135 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7485__A2 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5448_ _2095_ mod.Data_Mem.F_M.MRAM\[798\]\[0\] _2096_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_133_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4299__A2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout100 net101 net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_8167_ mod.Data_Mem.F_M.out_data\[77\] net29 net267 mod.Arithmetic.I_out\[77\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout111 net112 net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5379_ mod.Data_Mem.F_M.MRAM\[791\]\[7\] mod.Data_Mem.F_M.MRAM\[788\]\[7\] mod.Data_Mem.F_M.MRAM\[789\]\[7\]
+ mod.Data_Mem.F_M.MRAM\[790\]\[7\] _1915_ _1917_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xfanout122 net123 net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout133 net134 net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7118_ _3507_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout144 net146 net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout155 net159 net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_8098_ mod.Data_Mem.F_M.out_data\[8\] net55 net345 mod.Arithmetic.CN.I_in\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout166 net169 net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5248__A1 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout177 net178 net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6445__B1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5099__I1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout188 net189 net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6445__C2 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7049_ _3471_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout199 net200 net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_41_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5343__S1 _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5799__A2 _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6436__C _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__I0 mod.Data_Mem.F_M.MRAM\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5971__A2 mod.Data_Mem.F_M.MRAM\[773\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__C _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6359__S0 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5582__I _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5326__I2 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8115__CLK net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5031__S0 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5487__B2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__I mod.Arithmetic.CN.I_in\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6039__I0 mod.Data_Mem.F_M.MRAM\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4462__A2 _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4214__A2 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout337_I net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4750_ _1374_ _1378_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7539__I0 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3973__A1 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ _1226_ _0995_ _1232_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6420_ _1762_ _3025_ _3028_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5714__A2 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5706__B _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6351_ _2881_ _2960_ _2961_ _2879_ _1727_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5302_ mod.Data_Mem.F_M.MRAM\[5\]\[5\] mod.Data_Mem.F_M.MRAM\[4\]\[5\] _1570_ _1966_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6282_ _1607_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5478__A1 _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8021_ _0230_ net109 mod.Data_Mem.F_M.MRAM\[15\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5233_ _1888_ _1897_ _1635_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5164_ _1661_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6537__B _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4115_ mod.Arithmetic.ACTI.x\[5\] _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4046_ _0716_ _0718_ _0720_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__A1 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7778__I0 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7805_ mod.Data_Mem.F_M.MRAM\[7\]\[2\] _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5667__I _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5997_ _2524_ _2613_ _2615_ _2525_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5253__I1 mod.Data_Mem.F_M.MRAM\[788\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7736_ mod.Data_Mem.F_M.MRAM\[795\]\[4\] _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4948_ _1564_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5953__A2 mod.Data_Mem.F_M.MRAM\[21\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7667_ _3827_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ mod.Data_Mem.F_M.MRAM\[6\]\[0\] _1544_ _1547_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _3199_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7598_ _1686_ _3789_ _3790_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5705__A2 mod.Data_Mem.F_M.MRAM\[797\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6549_ _3083_ _3139_ _3141_ _3148_ _3151_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_106_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5335__C _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8219_ _0320_ net299 mod.Data_Mem.F_M.MRAM\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4947__S _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8508__573 net573 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__B1 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__C2 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5316__S1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7630__A2 _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5244__I1 mod.Data_Mem.F_M.MRAM\[768\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A2 mod.Data_Mem.F_M.MRAM\[14\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7146__A1 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7792__I _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4380__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4132__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5880__A1 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7032__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A1 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6871__I mod.Data_Mem.F_M.MRAM\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5920_ _2540_ mod.Data_Mem.F_M.MRAM\[773\]\[4\] _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5851_ mod.Data_Mem.F_M.MRAM\[4\]\[2\] mod.Data_Mem.F_M.MRAM\[5\]\[2\] mod.Data_Mem.F_M.MRAM\[20\]\[2\]
+ mod.Data_Mem.F_M.MRAM\[21\]\[2\] _1769_ _2104_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6188__A2 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _1454_ _1457_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4199__A1 mod.Arithmetic.CN.I_in\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8570_ _0074_ net349 mod.Data_Mem.F_M.out_data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5782_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5935__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7521_ _3741_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4733_ mod.Arithmetic.CN.I_in\[61\] _1366_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7452_ _3699_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4664_ mod.Arithmetic.CN.I_in\[38\] _1333_ _1334_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5699__A1 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6403_ _3008_ _2382_ _2377_ _2492_ _3011_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7383_ mod.Data_Mem.F_M.MRAM\[774\]\[0\] _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4595_ _1031_ _1263_ _1265_ _1266_ mod.P3.Res\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6334_ _2887_ _2003_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8430__CLK net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _2701_ _2684_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6112__A2 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__S _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8004_ _0213_ net232 mod.Data_Mem.F_M.MRAM\[13\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5216_ mod.Data_Mem.F_M.MRAM\[3\]\[4\] mod.Data_Mem.F_M.MRAM\[2\]\[4\] _1880_ _1881_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6196_ _1882_ _1753_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4674__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5871__A1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8580__CLK net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5871__B2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5147_ _1547_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5078_ _1602_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5623__A1 _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6781__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4029_ _0702_ mod.Arithmetic.I_out\[78\] _0703_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_38_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5397__I _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6179__A2 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__A2 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6974__I1 mod.Data_Mem.F_M.MRAM\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7719_ _3853_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7151__I1 mod.Data_Mem.F_M.MRAM\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4114__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__A2 mod.Arithmetic.CN.I_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8096__RN net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6691__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5614__B2 _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5100__I _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7027__I _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6342__A2 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout202_I net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4380_ _0617_ _0686_ _0688_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _2503_ mod.Data_Mem.F_M.MRAM\[4\]\[7\] _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_113_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5001_ _1589_ _1668_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4408__A2 _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5605__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6952_ _3386_ mod.Data_Mem.F_M.MRAM\[15\]\[0\] _3409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _2374_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4335__B mod.Arithmetic.ACTI.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6883_ mod.Data_Mem.F_M.MRAM\[4\]\[1\] _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5834_ _2454_ _2456_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5010__I _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6956__I1 mod.Data_Mem.F_M.MRAM\[15\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6030__B2 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ _2389_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8553_ _0057_ net342 mod.Data_Mem.F_M.out_data\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4592__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7504_ _3321_ _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4716_ _1325_ _1328_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8484_ _0580_ net101 mod.Data_Mem.F_M.MRAM\[798\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5696_ _2095_ mod.Data_Mem.F_M.MRAM\[797\]\[5\] _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7435_ mod.Data_Mem.F_M.MRAM\[777\]\[2\] _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _1313_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7366_ _3656_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4578_ _1241_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4895__A2 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6776__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6317_ _2883_ _2925_ _2928_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7297_ _3311_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5680__I _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A1 _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5144__I0 mod.Data_Mem.F_M.MRAM\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5613__C _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6248_ _2205_ _1628_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4647__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _2199_ _2675_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7601__S _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7597__A1 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8078__RN net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A2 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__I _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6947__I1 mod.Data_Mem.F_M.MRAM\[14\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6021__A1 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7048__S _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4335__A1 mod.Arithmetic.CN.I_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6686__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__A2 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7124__I1 mod.Data_Mem.F_M.MRAM\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A2 _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5835__A1 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_410 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7511__S _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_421 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_432 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_443 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_454 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_465 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_476 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8553__D _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_487 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4934__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_498 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout152_I net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A1 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6563__A2 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5765__I _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5550_ _1642_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4574__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4501_ _0684_ mod.Arithmetic.CN.I_in\[20\] _0613_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5481_ _2108_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6315__A2 _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7220_ _3252_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4326__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__I0 mod.Data_Mem.F_M.MRAM\[771\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4432_ _1018_ _1020_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7151_ _3527_ mod.Data_Mem.F_M.MRAM\[12\]\[1\] _3525_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4363_ _0863_ _0938_ _1027_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6102_ _2177_ _2717_ _2718_ _2710_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7082_ mod.Data_Mem.F_M.MRAM\[21\]\[4\] _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4294_ _0870_ _0966_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _2540_ mod.Data_Mem.F_M.MRAM\[773\]\[7\] _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5005__I mod.Data_Mem.F_M.src\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4049__C _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout65_I net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8499__CLK net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7220__I _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7984_ mod.Instr_Mem.instruction\[9\] net16 net218 mod.P1.instr_reg\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_54_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5054__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _3397_ mod.Data_Mem.F_M.MRAM\[14\]\[3\] _3391_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4801__A2 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6929__I1 mod.Data_Mem.F_M.MRAM\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6866_ _3355_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__A1 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6003__B2 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5817_ mod.Data_Mem.F_M.MRAM\[4\]\[1\] mod.Data_Mem.F_M.MRAM\[5\]\[1\] mod.Data_Mem.F_M.MRAM\[20\]\[1\]
+ mod.Data_Mem.F_M.MRAM\[21\]\[1\] _1923_ _2104_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_6797_ _3314_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6554__A2 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4565__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5748_ _2087_ _2058_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8536_ _0040_ net330 mod.Data_Mem.F_M.out_data\[32\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ _2210_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8467_ _0563_ net288 mod.Data_Mem.F_M.MRAM\[796\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4317__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7418_ _3682_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8398_ _0494_ net104 mod.Data_Mem.F_M.MRAM\[786\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7349_ _3620_ mod.Data_Mem.F_M.MRAM\[771\]\[7\] _3643_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7331__S _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__A2 mod.Data_Mem.F_M.MRAM\[768\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6490__A1 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__A1 _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__B2 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5585__I _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4703__B _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6545__A2 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7345__I1 mod.Data_Mem.F_M.MRAM\[771\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4859__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4929__I _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5284__A2 _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout367_I net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7040__I _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6233__A1 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4981_ _1510_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6720_ _3263_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4795__A1 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output6_I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7033__I0 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6651_ mod.Data_Mem.F_M.MRAM\[25\]\[5\] _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7584__I1 mod.Data_Mem.F_M.MRAM\[785\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ mod.Data_Mem.F_M.MRAM\[797\]\[5\] _2214_ _1750_ mod.Data_Mem.F_M.MRAM\[796\]\[5\]
+ _2237_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6582_ _3178_ _3179_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8321_ _0417_ net303 mod.Data_Mem.F_M.MRAM\[776\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5533_ _2163_ _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8252_ _0348_ net101 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6320__S _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _2109_ _2110_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8171__CLK net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7203_ _3537_ mod.Data_Mem.F_M.MRAM\[29\]\[6\] _3553_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4415_ _0986_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8183_ _0293_ net106 mod.Data_Mem.F_M.MRAM\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5395_ _2055_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5362__I3 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7134_ _3454_ mod.Data_Mem.F_M.MRAM\[19\]\[3\] _3513_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout304 net309 net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4346_ _0817_ _0923_ _0844_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_98_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout315 net318 net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout326 net391 net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout337 net338 net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout348 net350 net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__6847__I0 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7065_ _3479_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4277_ _0947_ _0949_ _0935_ _0950_ _0891_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
Xfanout359 net360 net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__7151__S _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6472__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5275__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6016_ _2498_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6472__B2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A1 mod.Data_Mem.F_M.MRAM\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7967_ _0193_ net144 mod.Data_Mem.F_M.MRAM\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4786__A1 mod.Arithmetic.CN.I_in\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6918_ _3259_ mod.Data_Mem.F_M.MRAM\[13\]\[7\] _3381_ _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7898_ _0124_ net383 mod.Data_Mem.F_M.MRAM\[27\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7024__I0 _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6849_ mod.Data_Mem.F_M.MRAM\[779\]\[0\] _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8519_ net566 net361 mod.Data_Mem.F_M.out_data\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7326__S _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5338__I0 mod.Data_Mem.F_M.MRAM\[771\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5889__I1 mod.Data_Mem.F_M.MRAM\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6169__C _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6463__A1 _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__B2 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7263__I0 mod.Data_Mem.F_M.MRAM\[31\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__I0 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4241__A3 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8194__CLK net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout115_I net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5264__B _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4200_ _0615_ _0873_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5180_ mod.Data_Mem.F_M.MRAM\[772\]\[3\] _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4131_ _0653_ _0676_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7246__A3 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4062_ _0731_ _0733_ _0736_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_95_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6206__A1 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__I0 mod.Data_Mem.F_M.MRAM\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7821_ _3910_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5965__B1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4964_ _1629_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7752_ _3309_ mod.Data_Mem.F_M.MRAM\[796\]\[3\] _3867_ _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6703_ net8 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8537__CLK net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7683_ _3835_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4895_ _1495_ _1505_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6634_ _3207_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5193__A1 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6565_ _3016_ _3163_ _3165_ _3166_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8304_ _0400_ net160 mod.Data_Mem.F_M.MRAM\[774\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5516_ _1682_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6496_ _3098_ _3099_ _3100_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8235_ _0331_ net213 mod.Data_Mem.F_M.MRAM\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6985__S _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5447_ _1908_ mod.Data_Mem.F_M.MRAM\[799\]\[0\] _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5496__A2 mod.Data_Mem.F_M.MRAM\[798\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout101 net103 net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_8166_ mod.Data_Mem.F_M.out_data\[76\] net28 net266 mod.Arithmetic.I_out\[76\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5378_ _1872_ _2039_ _1863_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xfanout112 net113 net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout123 net124 net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7117_ _3456_ mod.Data_Mem.F_M.MRAM\[3\]\[4\] _3506_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout134 net135 net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4329_ _0914_ _0920_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8097_ mod.Data_Mem.F_M.out_data\[7\] net26 net246 mod.Arithmetic.ACTI.x\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout145 net146 net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout156 net157 net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_113_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout167 net169 net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6445__A1 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7493__I0 _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7048_ _3454_ mod.Data_Mem.F_M.MRAM\[1\]\[3\] _3469_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout178 net216 net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_86_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6445__B2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout189 net200 net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8067__CLK net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__I1 mod.Data_Mem.F_M.MRAM\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4059__I0 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A2 _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5708__B1 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A1 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7056__S _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6359__S1 _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6133__B1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5326__I3 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5487__A2 _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5892__C1 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6694__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6436__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6039__I1 mod.Data_Mem.F_M.MRAM\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4462__A3 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8561__D _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7539__I1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5974__S _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout232_I net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3973__A2 mod.Arithmetic.CN.I_in\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4680_ _1228_ _1231_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5175__A1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6869__I mod.Data_Mem.F_M.MRAM\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6350_ _1992_ _1993_ _2895_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5301_ mod.Data_Mem.F_M.MRAM\[15\]\[5\] _1934_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4389__I mod.Arithmetic.CN.I_in\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6281_ mod.Data_Mem.F_M.MRAM\[789\]\[4\] mod.Data_Mem.F_M.MRAM\[791\]\[4\] mod.Data_Mem.F_M.MRAM\[790\]\[4\]
+ mod.Data_Mem.F_M.MRAM\[788\]\[4\] _2167_ _2376_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__6124__B1 _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5478__A2 _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8020_ _0229_ net109 mod.Data_Mem.F_M.MRAM\[15\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6675__A1 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5232_ _1891_ _1893_ _1894_ _1895_ _1896_ _1666_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_130_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4150__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5163_ _1662_ _1828_ _1664_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5214__S _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6427__A1 _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4114_ _0738_ _0784_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5094_ _1674_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4045_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5013__I _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5650__A2 _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6553__B _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7778__I1 mod.Data_Mem.F_M.MRAM\[797\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4852__I mod.Data_Mem.F_M.src\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7804_ _3900_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7927__CLK net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _2056_ mod.Data_Mem.F_M.MRAM\[772\]\[6\] _2614_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__I2 mod.Data_Mem.F_M.MRAM\[789\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7735_ _3861_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4947_ mod.Data_Mem.F_M.MRAM\[785\]\[0\] mod.Data_Mem.F_M.MRAM\[784\]\[0\] _1615_
+ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7666_ mod.Data_Mem.F_M.MRAM\[791\]\[1\] _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4878_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6617_ mod.Data_Mem.F_M.MRAM\[24\]\[4\] _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7597_ _3610_ _3789_ _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5616__C _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6548_ _1491_ _3150_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6479_ _2464_ mod.Data_Mem.F_M.MRAM\[769\]\[3\] _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8218_ _0319_ net81 mod.Data_Mem.F_M.MRAM\[22\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8149_ mod.Data_Mem.F_M.out_data\[59\] net57 net354 mod.Arithmetic.CN.I_in\[59\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__6418__A1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7466__I0 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5351__C _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6418__B2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7218__I0 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7769__I1 mod.Data_Mem.F_M.MRAM\[797\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5157__A1 _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4904__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5952__I0 mod.Data_Mem.F_M.MRAM\[16\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4380__A2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4002__I mod.Arithmetic.ACTI.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8556__D _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7313__I _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6409__A1 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5880__A2 _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout182_I net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__I0 _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5632__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _2372_ _2463_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _1459_ _1463_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_61_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4199__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _1490_ _2116_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7520_ _3645_ mod.Data_Mem.F_M.MRAM\[782\]\[5\] _3739_ _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4732_ _1400_ _1384_ _1401_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5148__A1 mod.Data_Mem.F_M.MRAM\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7451_ mod.Data_Mem.F_M.MRAM\[778\]\[2\] _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5148__B2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4663_ mod.Arithmetic.CN.I_in\[38\] _1333_ _1252_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5699__A2 _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _2414_ _3009_ _3010_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_128_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4594_ _0792_ _0857_ _0628_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7382_ _3664_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6333_ _1582_ _2002_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5008__I _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _1891_ _1893_ _1746_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_fanout95_I net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__B1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8003_ _0212_ net232 mod.Data_Mem.F_M.MRAM\[13\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5215_ _1873_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5320__A1 _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6195_ _2582_ mod.Data_Mem.F_M.MRAM\[22\]\[2\] mod.Data_Mem.F_M.MRAM\[23\]\[2\] _2753_
+ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ mod.Data_Mem.F_M.MRAM\[5\]\[3\] mod.Data_Mem.F_M.MRAM\[4\]\[3\] _1611_ _1812_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5871__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5077_ mod.Data_Mem.F_M.MRAM\[17\]\[2\] mod.Data_Mem.F_M.MRAM\[16\]\[2\] _1658_ _1744_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5623__A2 _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4028_ _0702_ mod.Arithmetic.I_out\[78\] _0684_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7620__I0 _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8105__CLK net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5979_ _2399_ _2597_ _2598_ _2396_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7718_ mod.Data_Mem.F_M.MRAM\[794\]\[3\] _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7649_ _3818_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__S _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__A3 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5311__A1 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5614__A2 mod.Data_Mem.F_M.MRAM\[799\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7509__S _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5925__I0 mod.Data_Mem.F_M.MRAM\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7244__S _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6350__I0 _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5000_ mod.Data_Mem.F_M.MRAM\[21\]\[1\] mod.Data_Mem.F_M.MRAM\[20\]\[1\] _1639_ _1668_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6951_ _3408_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_54_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5498__I _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _1728_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6882_ _3363_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4335__C _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5833_ _2410_ _1793_ _2455_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6030__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8552_ _0056_ net256 mod.Data_Mem.F_M.out_data\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5764_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7503_ _3730_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4715_ _1347_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8483_ _0579_ net256 mod.Data_Mem.F_M.MRAM\[798\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5695_ _2319_ _2321_ _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7434_ _3690_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5916__I0 mod.Data_Mem.F_M.MRAM\[770\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4646_ _1061_ _1314_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_116_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5541__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7365_ mod.Data_Mem.F_M.MRAM\[772\]\[7\] _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4577_ _1242_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7154__S _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _2713_ _2926_ _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7296_ _1855_ _3609_ _3614_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7294__A1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6097__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__I1 mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6247_ _1865_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6178_ _2067_ _2788_ _2792_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6792__I _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5129_ _1763_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7597__A2 _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A2 _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6460__C _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A3 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_400 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_411 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_422 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_433 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_444 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_455 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__S _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_466 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_477 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5599__A1 mod.Data_Mem.F_M.MRAM\[29\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_488 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5599__B2 mod.Data_Mem.F_M.MRAM\[28\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_499 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6012__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout145_I net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4023__A1 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5071__I0 mod.Data_Mem.F_M.MRAM\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4574__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8570__CLK net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7038__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout312_I net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4500_ _1170_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5480_ mod.Data_Mem.F_M.MRAM\[30\]\[3\] mod.Data_Mem.F_M.MRAM\[31\]\[3\] _1787_ _2126_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4431_ _0828_ _1018_ _1020_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4326__A2 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__I1 mod.Data_Mem.F_M.MRAM\[770\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7150_ _3239_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4362_ _0945_ _1026_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6101_ _1740_ _1571_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7081_ _3487_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4293_ _0880_ _0881_ _0872_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ mod.Data_Mem.F_M.MRAM\[770\]\[7\] mod.Data_Mem.F_M.MRAM\[771\]\[7\] _2490_
+ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout58_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7983_ mod.Instr_Mem.instruction\[8\] net34 net263 mod.P1.instr_reg\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_81_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6934_ _3245_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ mod.Data_Mem.F_M.MRAM\[6\]\[0\] _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4860__I _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _2088_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6796_ mod.Data_Mem.F_M.MRAM\[799\]\[4\] _3312_ _3313_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8535_ _0039_ net254 mod.Data_Mem.F_M.out_data\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5747_ _2371_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7991__RN net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8466_ _0562_ net292 mod.Data_Mem.F_M.MRAM\[796\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5678_ _2301_ _2307_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7417_ mod.Data_Mem.F_M.MRAM\[776\]\[1\] _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4629_ _1185_ _1093_ _1184_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8511__570 net570 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_8397_ _0493_ net105 mod.Data_Mem.F_M.MRAM\[786\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7348_ _3647_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ mod.Data_Mem.F_M.MRAM\[5\]\[7\] _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5640__B _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8443__CLK net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__A2 mod.Data_Mem.F_M.MRAM\[783\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8593__CLK net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5866__I _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4005__A1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4703__C mod.Arithmetic.ACTI.x\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A2 mod.Arithmetic.CN.I_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7982__RN net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5505__A1 _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput3 net3 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7522__S _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4945__I _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4492__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5977__S _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout262_I net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4980_ _1647_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7033__I1 mod.Data_Mem.F_M.MRAM\[18\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _3215_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7960__CLK net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__A3 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5601_ _1708_ _2236_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4547__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _3175_ _3176_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8320_ _0416_ net375 mod.Data_Mem.F_M.MRAM\[776\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5532_ _2154_ _2164_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8251_ _0347_ net311 mod.Data_Mem.F_M.MRAM\[31\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ _2111_ _2060_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7202_ _3558_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4414_ _0992_ _1085_ _1086_ _1023_ _0988_ _0989_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
X_8182_ _0292_ net109 mod.Data_Mem.F_M.MRAM\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5394_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7133_ _3516_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout305 net307 net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4345_ _0649_ _1017_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout316 net318 net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout327 net328 net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6847__I1 mod.Data_Mem.F_M.MRAM\[769\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout338 net353 net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7064_ mod.Data_Mem.F_M.MRAM\[20\]\[3\] _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4276_ _0904_ _0934_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xfanout349 net351 net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_101_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8150__RN net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6015_ _2579_ mod.Data_Mem.F_M.MRAM\[5\]\[6\] _2633_ _2089_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6048__S _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6224__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7966_ _0192_ net164 mod.Data_Mem.F_M.MRAM\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4235__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__I0 mod.Data_Mem.F_M.MRAM\[785\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ _3384_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7897_ _0123_ net193 mod.Data_Mem.F_M.MRAM\[27\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5686__I _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7024__I1 mod.Data_Mem.F_M.MRAM\[18\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6848_ _3346_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A2 mod.Arithmetic.CN.I_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ mod.Data_Mem.F_M.MRAM\[799\]\[0\] _3293_ _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6783__I0 mod.Data_Mem.F_M.MRAM\[799\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7607__S _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8518_ net567 net362 mod.Data_Mem.F_M.out_data\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8449_ _0545_ net376 mod.Data_Mem.F_M.MRAM\[794\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5338__I1 mod.Data_Mem.F_M.MRAM\[770\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5889__I2 mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5354__C _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6160__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7342__S _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5370__B _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__A2 _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8141__RN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6215__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7263__I1 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7983__CLK net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7015__I1 mod.Data_Mem.F_M.MRAM\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8339__CLK net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8559__D _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5037__S _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout108_I net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__S _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4130_ _0629_ _0677_ _0806_ mod.P3.Res\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4061_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6206__A2 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7254__I1 _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7820_ _3907_ _3908_ _3909_ _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_64_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7751_ _3870_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4963_ _1631_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5965__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5965__B2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6702_ _3251_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7682_ mod.Data_Mem.F_M.MRAM\[792\]\[1\] _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4894_ _1551_ _1557_ _1562_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6633_ mod.Data_Mem.F_M.MRAM\[26\]\[4\] _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8199__RN net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6564_ _2492_ _2649_ _2650_ _3008_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8303_ _0399_ net83 mod.Data_Mem.F_M.MRAM\[773\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5515_ _1526_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ _2500_ mod.Data_Mem.F_M.MRAM\[2\]\[4\] _2550_ _2560_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6130__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8234_ _0330_ net300 mod.Data_Mem.F_M.MRAM\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5446_ _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6142__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ mod.Data_Mem.F_M.out_data\[75\] net28 net266 mod.Arithmetic.I_out\[75\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5377_ _2035_ _2036_ _2037_ _2038_ _1911_ _1591_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xfanout102 net103 net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout113 net131 net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7116_ _3500_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xfanout124 net129 net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout135 net136 net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4328_ _1000_ _1001_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8096_ mod.Data_Mem.F_M.out_data\[6\] net26 net266 mod.Arithmetic.ACTI.x\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout146 net153 net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout157 net159 net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout168 net169 net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_87_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6445__A2 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ _3470_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7493__I1 mod.Data_Mem.F_M.MRAM\[781\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout179 net181 net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4259_ _0908_ _0927_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_80_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7949_ _0175_ net88 mod.Data_Mem.F_M.MRAM\[789\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5956__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__A1 _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5708__B2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7337__S _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A1 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6381__B2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4392__B1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7136__I _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6133__A1 mod.Data_Mem.F_M.MRAM\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6133__B2 mod.Data_Mem.F_M.MRAM\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__B1 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5892__C2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6436__A2 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout225_I net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6372__A1 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5300_ _1632_ _1951_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6124__A1 mod.Data_Mem.F_M.MRAM\[781\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6280_ _2878_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6124__B2 mod.Data_Mem.F_M.MRAM\[780\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6675__A2 mod.Data_Mem.F_M.dest\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5231_ _1601_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4686__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ mod.Data_Mem.F_M.MRAM\[787\]\[3\] mod.Data_Mem.F_M.MRAM\[786\]\[3\] _1615_
+ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__A2 mod.Data_Mem.F_M.MRAM\[769\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8105__RN net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7624__A1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4113_ _0736_ _0784_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5093_ _1756_ _1759_ _1598_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4044_ mod.Arithmetic.CN.I_in\[10\] _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8504__CLK net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__S _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout40_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7803_ mod.Data_Mem.F_M.MRAM\[7\]\[1\] _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _2418_ mod.Data_Mem.F_M.MRAM\[773\]\[6\] _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7734_ mod.Data_Mem.F_M.MRAM\[795\]\[3\] _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4946_ _1603_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7665_ _3826_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4877_ _1545_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7157__S _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6616_ _3198_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6363__A1 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7596_ _3786_ _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6996__S _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6547_ _3049_ _3149_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6115__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7163__I0 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _2351_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8217_ _0318_ net78 mod.Data_Mem.F_M.MRAM\[22\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6795__I _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5429_ _2081_ _2083_ _2070_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8034__CLK net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8148_ mod.Data_Mem.F_M.out_data\[58\] net55 net335 mod.Arithmetic.CN.I_in\[58\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_0_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6418__A2 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7466__I1 mod.Data_Mem.F_M.MRAM\[780\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8079_ mod.P3.Res\[7\] net26 net245 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_75_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7620__S _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__I0 mod.Data_Mem.F_M.MRAM\[798\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8184__CLK net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7218__I1 mod.Data_Mem.F_M.MRAM\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5157__A2 _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4904__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6106__A1 _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7154__I0 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4380__A3 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5315__S _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5542__C _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__A2 mod.Data_Mem.F_M.MRAM\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8572__D _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7209__I1 mod.Data_Mem.F_M.MRAM\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4953__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout175_I net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__I0 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _1464_ _1466_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA_fanout342_I net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4199__A3 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5780_ _2372_ _2386_ _2404_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _1347_ _1385_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5784__I _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7450_ _3698_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5148__A2 _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6345__A1 _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4662_ _1090_ _1331_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6401_ _2207_ mod.Data_Mem.F_M.MRAM\[781\]\[0\] _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7381_ mod.Data_Mem.F_M.MRAM\[773\]\[7\] _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _0792_ _0805_ _0859_ _1264_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6332_ _2864_ _2943_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6263_ _2867_ _2875_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4659__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8002_ _0211_ net305 mod.Data_Mem.F_M.MRAM\[13\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4659__B2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5214_ mod.Data_Mem.F_M.MRAM\[1\]\[4\] mod.Data_Mem.F_M.MRAM\[0\]\[4\] _1878_ _1879_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6194_ _2757_ _2807_ _2808_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5145_ mod.Data_Mem.F_M.MRAM\[22\]\[3\] _1600_ _1614_ _1810_ _1508_ _1811_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_57_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5024__I _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5076_ _1735_ _1736_ _1739_ _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5959__I _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__A1 mod.Data_Mem.F_M.MRAM\[22\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4027_ mod.Arithmetic.I_out\[77\] _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5895__S _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5978_ mod.Data_Mem.F_M.MRAM\[784\]\[5\] mod.Data_Mem.F_M.MRAM\[785\]\[5\] _2224_
+ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7717_ _3852_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4929_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6336__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7648_ mod.Data_Mem.F_M.MRAM\[790\]\[0\] _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7579_ _3777_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7615__S _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7836__A1 _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3942__I _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5075__A1 _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6590__A4 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6327__A1 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4889__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4013__I mod.Arithmetic.CN.I_in\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4948__I _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7917__CLK net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout292_I net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6950_ _3235_ _3407_ _3374_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5901_ _2074_ _2509_ _2522_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6881_ mod.Data_Mem.F_M.MRAM\[4\]\[0\] _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _2304_ mod.Data_Mem.F_M.MRAM\[787\]\[2\] _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6566__A1 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8551_ _0055_ net251 mod.Data_Mem.F_M.out_data\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5763_ _1594_ _1495_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7502_ _3729_ mod.Data_Mem.F_M.MRAM\[781\]\[6\] _3726_ _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4714_ _1349_ _1384_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8482_ _0578_ net341 mod.Data_Mem.F_M.MRAM\[798\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5694_ _2115_ _2141_ _2143_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7433_ mod.Data_Mem.F_M.MRAM\[777\]\[1\] _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4645_ _1063_ _1178_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5916__I1 mod.Data_Mem.F_M.MRAM\[771\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7364_ _3655_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4576_ _1243_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6315_ _2889_ _1958_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7295_ _3555_ _3606_ _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7294__A2 _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _2846_ _2853_ _2859_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6341__I1 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6177_ _2680_ _2791_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5128_ _1791_ mod.Data_Mem.F_M.MRAM\[787\]\[2\] _1794_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5057__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _1673_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5852__I0 mod.Data_Mem.F_M.MRAM\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6557__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3937__I _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7345__S _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5532__A2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4638__A4 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_401 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_412 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_423 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_434 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5048__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_445 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_456 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_467 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_63_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_478 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_489 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6340__S0 _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4008__I _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__I1 mod.Data_Mem.F_M.MRAM\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5267__C _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout138_I net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4879__S _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout305_I net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4430_ _1089_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4361_ _0787_ _0856_ _0858_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6100_ _2705_ mod.Data_Mem.F_M.MRAM\[774\]\[0\] mod.Data_Mem.F_M.MRAM\[775\]\[0\]
+ _2158_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7080_ mod.Data_Mem.F_M.MRAM\[21\]\[3\] _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7520__I0 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4292_ _0872_ _0880_ _0881_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5287__A1 _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ mod.Data_Mem.F_M.MRAM\[782\]\[7\] mod.Data_Mem.F_M.MRAM\[783\]\[7\] _2571_
+ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6893__I mod.Data_Mem.F_M.MRAM\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7982_ mod.Instr_Mem.instruction\[7\] net25 net263 mod.P1.instr_reg\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8245__CLK net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6933_ _3396_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6864_ _3354_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__A1 _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7587__I0 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5815_ _2409_ _2424_ _2438_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6795_ _3299_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8534_ _0038_ net253 mod.Data_Mem.F_M.out_data\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5746_ _2370_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7339__I0 _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8465_ _0561_ net291 mod.Data_Mem.F_M.MRAM\[796\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5677_ _2302_ _2306_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7416_ _3681_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4628_ _1185_ _1093_ _1184_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8396_ _0492_ net104 mod.Data_Mem.F_M.MRAM\[786\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5514__A2 _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7347_ _3618_ mod.Data_Mem.F_M.MRAM\[771\]\[6\] _3643_ _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4559_ _1229_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7511__I0 _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7278_ _3601_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5278__A1 _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6229_ _1805_ _1832_ _2842_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__I0 mod.Data_Mem.F_M.MRAM\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__A1 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7578__I0 _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4005__A2 mod.Arithmetic.I_out\[79\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6389__S0 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5505__A2 mod.Data_Mem.F_M.MRAM\[798\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7750__I0 _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8118__CLK net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput4 net4 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7502__I0 _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5323__S _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout255_I net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__C _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5600_ _2229_ mod.Data_Mem.F_M.MRAM\[799\]\[5\] mod.Data_Mem.F_M.MRAM\[798\]\[5\]
+ _1816_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_34_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6580_ mod.I_addr\[4\] _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4547__A3 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5531_ mod.Data_Mem.F_M.MRAM\[797\]\[0\] _1731_ _2171_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8250_ _0346_ net341 mod.Data_Mem.F_M.MRAM\[31\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5462_ _1806_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7201_ _3508_ mod.Data_Mem.F_M.MRAM\[29\]\[5\] _3553_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4413_ _1002_ _1022_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8181_ _0291_ net206 mod.Data_Mem.F_M.MRAM\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5393_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7132_ _3452_ mod.Data_Mem.F_M.MRAM\[19\]\[2\] _3513_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4344_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout306 net307 net306 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout317 net318 net317 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6457__B1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout328 net329 net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout339 net343 net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_7063_ _3478_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4275_ _0868_ _0888_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6556__C _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout70_I net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6014_ _2632_ mod.Data_Mem.F_M.MRAM\[4\]\[6\] _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_101_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7965_ _0191_ net369 mod.Data_Mem.F_M.MRAM\[779\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4235__A2 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5283__I1 mod.Data_Mem.F_M.MRAM\[784\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6916_ _3256_ mod.Data_Mem.F_M.MRAM\[13\]\[6\] _3381_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7896_ _0122_ net369 mod.Data_Mem.F_M.MRAM\[27\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5983__A2 _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6847_ _3259_ mod.Data_Mem.F_M.MRAM\[769\]\[7\] _3336_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _3299_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6783__I1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6798__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5729_ mod.Data_Mem.F_M.MRAM\[16\]\[0\] mod.Data_Mem.F_M.MRAM\[17\]\[0\] _2353_ _2354_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8517_ net568 net362 mod.Data_Mem.F_M.out_data\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8448_ _0544_ net372 mod.Data_Mem.F_M.MRAM\[794\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5499__A1 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5889__I3 mod.Data_Mem.F_M.MRAM\[21\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8379_ _0475_ net180 mod.Data_Mem.F_M.MRAM\[784\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5207__I _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6160__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4171__A1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8410__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5671__A1 _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4982__S _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__I0 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6215__A3 mod.Data_Mem.F_M.MRAM\[20\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5877__I _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3985__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8090__CLK net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__B _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8575__D _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4060_ mod.Arithmetic.CN.I_in\[13\] _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4217__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ _1491_ _1499_ _1563_ _1626_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_7750_ _3749_ mod.Data_Mem.F_M.MRAM\[796\]\[2\] _3867_ _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5965__A2 _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6701_ _3249_ mod.Data_Mem.F_M.MRAM\[28\]\[4\] _3250_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__3976__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7681_ _3834_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4893_ mod.Data_Mem.F_M.MRAM\[15\]\[0\] _1536_ mod.Data_Mem.F_M.MRAM\[31\]\[0\] _1561_
+ _1556_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ _3206_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5717__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ mod.Data_Mem.F_M.MRAM\[780\]\[7\] _1680_ _2559_ _3164_ _2617_ _3165_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5228__S _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6411__I _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8302_ _0398_ net86 mod.Data_Mem.F_M.MRAM\[773\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5514_ _2154_ _2091_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6494_ _3084_ mod.Data_Mem.F_M.MRAM\[0\]\[4\] _2101_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8233_ _0329_ net204 mod.Data_Mem.F_M.MRAM\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5445_ _1522_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6142__A2 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5027__I _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4153__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8164_ mod.Data_Mem.F_M.out_data\[74\] net31 net270 mod.Arithmetic.I_out\[74\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5376_ mod.Data_Mem.F_M.MRAM\[775\]\[7\] mod.Data_Mem.F_M.MRAM\[774\]\[7\] _1831_
+ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout103 net113 net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7115_ _3505_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8583__CLK net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__I _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout114 net115 net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4327_ _0993_ _0999_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout125 net128 net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_8095_ mod.Data_Mem.F_M.out_data\[5\] net51 net282 mod.Arithmetic.ACTI.x\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout136 net137 net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout147 net148 net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout158 net177 net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _3452_ mod.Data_Mem.F_M.MRAM\[1\]\[2\] _3469_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout169 net175 net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4258_ _0929_ _0931_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_86_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4456__A2 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5653__A1 _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ _0808_ _0822_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5697__I _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7948_ _0174_ net85 mod.Data_Mem.F_M.MRAM\[789\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7879_ _0105_ net317 mod.Data_Mem.F_M.MRAM\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7618__S _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5708__A2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6381__A2 _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3945__I _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4392__B2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6133__A2 _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4144__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__A1 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5892__B2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7950__CLK net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5644__A1 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6692__I0 _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6991__I _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8306__CLK net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5247__I1 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7528__S _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4016__I _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6372__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7327__I _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout120_I net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4383__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout218_I net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6124__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7263__S _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ mod.Data_Mem.F_M.MRAM\[17\]\[4\] mod.Data_Mem.F_M.MRAM\[16\]\[4\] _1718_ _1895_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5883__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ _1657_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4112_ _0777_ _0783_ _0786_ _0787_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7624__A2 _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _1758_ mod.Data_Mem.F_M.MRAM\[31\]\[2\] _1724_ mod.Data_Mem.F_M.MRAM\[15\]\[2\]
+ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5635__A1 _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _0693_ _0689_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4635__B _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7802_ _3899_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ _2611_ mod.Data_Mem.F_M.MRAM\[782\]\[6\] _2612_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6060__A1 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout33_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7733_ _3860_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4945_ _1601_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A2 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4876_ _1503_ _1504_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7664_ mod.Data_Mem.F_M.MRAM\[791\]\[0\] _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6615_ mod.Data_Mem.F_M.MRAM\[24\]\[3\] _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7595_ _3788_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7237__I _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__A2 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6141__I _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6546_ _3047_ _2334_ _2488_ _2607_ _2608_ _2559_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6477_ _2693_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7163__I1 mod.Data_Mem.F_M.MRAM\[12\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7973__CLK net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8216_ _0317_ net89 mod.Data_Mem.F_M.MRAM\[22\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5428_ _2082_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4921__I0 mod.Data_Mem.F_M.MRAM\[769\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ mod.Data_Mem.F_M.MRAM\[3\]\[7\] mod.Data_Mem.F_M.MRAM\[2\]\[7\] _1876_ _2021_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8147_ mod.Data_Mem.F_M.out_data\[57\] net52 net334 mod.Arithmetic.CN.I_in\[57\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_99_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8078_ mod.P3.Res\[6\] net34 net262 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_82_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__I1 mod.Data_Mem.F_M.MRAM\[799\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7029_ _3458_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5229__I1 mod.Data_Mem.F_M.MRAM\[18\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4037__S _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6051__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__B1 _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4601__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7147__I _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6354__A2 _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6106__A2 mod.Data_Mem.F_M.MRAM\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7154__I1 mod.Data_Mem.F_M.MRAM\[12\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4117__A1 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A2 mod.Arithmetic.CN.I_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8099__RN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5617__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5617__B2 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5331__S _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6968__I1 mod.Data_Mem.F_M.MRAM\[15\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6042__A1 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout335_I net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4730_ _1349_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _0659_ mod.Arithmetic.CN.I_in\[35\] _1090_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6400_ _2705_ mod.Data_Mem.F_M.MRAM\[780\]\[0\] _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4356__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7380_ _3663_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5553__B1 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4592_ _0791_ _0801_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _2866_ _2934_ _2942_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_157_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4108__A1 _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6262_ _2869_ _2871_ _2872_ _2874_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8001_ _0210_ net297 mod.Data_Mem.F_M.MRAM\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5213_ _1584_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6193_ _2178_ _1744_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ mod.Data_Mem.F_M.MRAM\[21\]\[3\] mod.Data_Mem.F_M.MRAM\[20\]\[3\] _1809_ _1810_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5608__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ _1740_ _1741_ _1617_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5084__A2 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4026_ mod.Arithmetic.CN.I_in\[23\] _0683_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5040__I _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6033__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6584__A2 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5977_ mod.Data_Mem.F_M.MRAM\[786\]\[5\] mod.Data_Mem.F_M.MRAM\[787\]\[5\] _1515_
+ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7716_ mod.Data_Mem.F_M.MRAM\[794\]\[2\] _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4928_ _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7647_ _3817_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6336__A2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4859_ _1502_ _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5544__B1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7578_ _3765_ mod.Data_Mem.F_M.MRAM\[785\]\[3\] _3773_ _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6529_ _2523_ _3123_ _3132_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7836__A2 mod.I_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5847__A1 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8151__CLK net361 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__I _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6272__A1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A2 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5783__B1 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4338__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4889__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5125__I _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4510__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout285_I net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5900_ _2515_ _2521_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6880_ _3362_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6015__A1 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ _2107_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6566__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8024__CLK net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4577__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8550_ _0054_ net252 mod.Data_Mem.F_M.out_data\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5762_ _2373_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7501_ _3318_ _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ _1363_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5693_ _2320_ mod.Data_Mem.F_M.MRAM\[28\]\[5\] _2254_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8481_ _0577_ net294 mod.Data_Mem.F_M.MRAM\[798\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6318__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7432_ _3689_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5377__I0 _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4644_ mod.Arithmetic.CN.I_in\[30\] _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8174__CLK net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7363_ mod.Data_Mem.F_M.MRAM\[772\]\[6\] _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4575_ _1244_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6314_ _1638_ _1959_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7294_ _1775_ _3609_ _3613_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6245_ _2106_ _2217_ _2858_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4501__A1 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6176_ mod.Data_Mem.F_M.MRAM\[781\]\[2\] _1731_ _2195_ mod.Data_Mem.F_M.MRAM\[780\]\[2\]
+ _2790_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_69_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ _1792_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5058_ mod.Data_Mem.F_M.MRAM\[783\]\[1\] _1702_ _1725_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5852__I1 mod.Data_Mem.F_M.MRAM\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4009_ mod.Arithmetic.CN.I_in\[19\] _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6006__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7054__I0 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4280__A3 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6557__A2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4568__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A4 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7626__S _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5368__I0 mod.Data_Mem.F_M.MRAM\[17\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5654__B _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3953__I mod.Arithmetic.CN.I_in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__S _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4050__S _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4740__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6493__A1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_402 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_413 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_424 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7160__I _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_435 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_446 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6245__A1 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5048__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_457 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_468 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_479 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6340__S1 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6705__S _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5220__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8197__CLK net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5851__S0 _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4024__I mod.Arithmetic.CN.I_in\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7536__S _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5359__I0 mod.Data_Mem.F_M.MRAM\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8578__D _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4959__I _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout200_I net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ _0786_ _0801_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4291_ _0953_ _0955_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_98_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7520__I1 mod.Data_Mem.F_M.MRAM\[782\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6030_ _2524_ _2152_ _2525_ _2643_ _2647_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6484__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7070__I mod.Data_Mem.F_M.MRAM\[20\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__A1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7981_ _0207_ net81 mod.Data_Mem.F_M.MRAM\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6932_ _3395_ mod.Data_Mem.F_M.MRAM\[14\]\[2\] _3391_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4798__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7036__I0 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6863_ mod.Data_Mem.F_M.MRAM\[779\]\[7\] _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__A2 mod.Data_Mem.F_M.MRAM\[781\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6414__I _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5814_ _2425_ _2437_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6794_ _3311_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8533_ _0037_ net277 mod.Data_Mem.F_M.out_data\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5745_ _2104_ _2369_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7339__I1 mod.Data_Mem.F_M.MRAM\[771\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6350__S _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8464_ _0560_ net287 mod.Data_Mem.F_M.MRAM\[796\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5676_ _2085_ _2130_ _2303_ _2305_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_108_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7415_ mod.Data_Mem.F_M.MRAM\[776\]\[0\] _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4869__I _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4627_ _1294_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8395_ _0491_ net179 mod.Data_Mem.F_M.MRAM\[786\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7346_ _3646_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4558_ mod.Arithmetic.CN.I_in\[53\] _1114_ _1116_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7277_ mod.Data_Mem.F_M.MRAM\[5\]\[6\] _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4489_ _1048_ _1077_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7511__I1 mod.Data_Mem.F_M.MRAM\[782\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5278__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6475__A1 _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6228_ _2709_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6159_ _2774_ _1721_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6227__A1 _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__I1 mod.Data_Mem.F_M.MRAM\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5450__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5649__B _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7907__CLK net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__A2 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A4 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4961__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__S1 _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4713__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput5 net5 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7502__I1 mod.Data_Mem.F_M.MRAM\[781\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6218__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7018__I0 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout150_I net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout248_I net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _2165_ _2170_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4952__A1 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5461_ mod.Data_Mem.F_M.MRAM\[30\]\[0\] mod.Data_Mem.F_M.MRAM\[31\]\[0\] _1712_ _2110_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7200_ _3557_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8101__D mod.Data_Mem.F_M.out_data\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4412_ _1002_ _1022_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4704__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8180_ _0290_ net207 mod.Data_Mem.F_M.MRAM\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5392_ _1522_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5752__I0 mod.Data_Mem.F_M.MRAM\[782\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7131_ _3515_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4343_ mod.Arithmetic.CN.I_in\[59\] _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout307 net308 net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6457__A1 mod.Data_Mem.F_M.MRAM\[13\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8212__CLK net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout318 net319 net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6457__B2 mod.Data_Mem.F_M.MRAM\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7062_ mod.Data_Mem.F_M.MRAM\[20\]\[2\] _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4274_ _0946_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xfanout329 net333 net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_99_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6013_ _1763_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7257__I0 mod.Data_Mem.F_M.MRAM\[31\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout63_I net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7964_ _0190_ net167 mod.Data_Mem.F_M.MRAM\[779\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7009__I0 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4235__A3 mod.Arithmetic.CN.I_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6915_ _3383_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7895_ _0121_ net370 mod.Data_Mem.F_M.MRAM\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6846_ _3345_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5196__A1 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6777_ _3294_ _3296_ _3298_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3989_ _0664_ _0665_ mod.Arithmetic.CN.I_in\[64\] _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8516_ net569 net359 mod.Data_Mem.F_M.out_data\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5728_ _1512_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_164_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8447_ _0543_ net342 mod.Data_Mem.F_M.MRAM\[793\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5659_ _2289_ mod.Data_Mem.F_M.MRAM\[29\]\[2\] _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__A2 mod.Data_Mem.F_M.MRAM\[31\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8378_ _0474_ net316 mod.Data_Mem.F_M.MRAM\[784\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7329_ _3272_ _3296_ _3634_ _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4171__A2 mod.Arithmetic.ACTI.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6448__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__I _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5671__A2 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7248__I0 mod.Data_Mem.F_M.MRAM\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__I1 mod.Data_Mem.F_M.MRAM\[798\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A2 mod.Arithmetic.CN.I_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8518__567 net567 vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__5187__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8235__CLK net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4162__A2 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7487__I0 _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8385__CLK net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5111__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout198_I net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6298__S0 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout365_I net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4961_ _1490_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _3236_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_33_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7680_ mod.Data_Mem.F_M.MRAM\[792\]\[0\] _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output4_I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4892_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6631_ mod.Data_Mem.F_M.MRAM\[26\]\[3\] _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4225__I0 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6562_ _2391_ mod.Data_Mem.F_M.MRAM\[768\]\[7\] _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8301_ _0397_ net142 mod.Data_Mem.F_M.MRAM\[773\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5513_ _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6493_ _2611_ mod.Data_Mem.F_M.MRAM\[1\]\[4\] _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8232_ _0328_ net296 mod.Data_Mem.F_M.MRAM\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5444_ _2089_ _2092_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8163_ mod.Data_Mem.F_M.out_data\[73\] net29 net270 mod.Arithmetic.I_out\[73\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__5350__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4153__A2 mod.Arithmetic.CN.I_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ mod.Data_Mem.F_M.MRAM\[773\]\[7\] mod.Data_Mem.F_M.MRAM\[772\]\[7\] _1908_
+ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5244__S _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7114_ _3454_ mod.Data_Mem.F_M.MRAM\[3\]\[3\] _3501_ _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xfanout104 net108 net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__7478__I0 _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout115 net117 net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4326_ _0993_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout126 net128 net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_8094_ mod.Data_Mem.F_M.out_data\[4\] net28 net268 mod.Arithmetic.ACTI.x\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
Xfanout137 net217 net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout148 net152 net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout159 net177 net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_7045_ _3465_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_59_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4257_ _0828_ _0929_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5043__I _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A2 mod.Data_Mem.F_M.MRAM\[797\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4188_ _0807_ _0854_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8108__CLK net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7947_ _0173_ net138 mod.Data_Mem.F_M.MRAM\[789\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7878_ _0104_ net372 mod.Data_Mem.F_M.MRAM\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6829_ _3334_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_23_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4144__A2 mod.Arithmetic.CN.I_in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5154__S _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__A2 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6692__I1 mod.Data_Mem.F_M.MRAM\[28\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5888__I _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__I2 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5947__A3 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6713__S _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5329__S _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4383__A2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7544__S _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4032__I _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout113_I net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4967__I _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ mod.Data_Mem.F_M.MRAM\[785\]\[3\] mod.Data_Mem.F_M.MRAM\[784\]\[3\] _1769_
+ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4111_ _0782_ _0780_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5091_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4042_ _0708_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4635__C _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7801_ mod.Data_Mem.F_M.MRAM\[7\]\[0\] _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5399__A1 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5993_ _1937_ mod.Data_Mem.F_M.MRAM\[783\]\[6\] _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_91_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7732_ mod.Data_Mem.F_M.MRAM\[795\]\[2\] _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4944_ _1608_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4071__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout26_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7663_ _3825_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4875_ mod.Data_Mem.F_M.MRAM\[5\]\[0\] mod.Data_Mem.F_M.MRAM\[4\]\[0\] _1543_ _1544_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6899__A1 mod.Data_Mem.F_M.dest\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6614_ _3197_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7594_ _3771_ mod.Data_Mem.F_M.MRAM\[786\]\[0\] _3787_ _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6545_ _2603_ _2619_ _3144_ _2204_ _3147_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4374__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _1676_ _3079_ _3081_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8215_ _0316_ net72 mod.Data_Mem.F_M.MRAM\[22\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4877__I _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _1554_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8146_ mod.Data_Mem.F_M.out_data\[56\] net67 net344 mod.Arithmetic.CN.I_in\[56\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ mod.Data_Mem.F_M.MRAM\[1\]\[7\] mod.Data_Mem.F_M.MRAM\[0\]\[7\] _1892_ _2020_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4309_ _0634_ mod.Arithmetic.CN.I_in\[43\] _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8077_ mod.P3.Res\[5\] net26 net264 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_5289_ mod.Data_Mem.F_M.MRAM\[775\]\[5\] mod.Data_Mem.F_M.MRAM\[774\]\[5\] _1585_
+ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7028_ _3456_ mod.Data_Mem.F_M.MRAM\[18\]\[4\] _3457_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8080__CLK net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4062__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4062__B2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3956__I _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5562__A1 _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5411__I _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7539__S _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8573__CLK net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout230_I net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ mod.Arithmetic.CN.I_in\[37\] _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_fanout328_I net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5553__A1 mod.Data_Mem.F_M.MRAM\[797\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _1261_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _2865_ _2941_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5305__A1 _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6261_ _2873_ _1879_ _2767_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8000_ _0209_ net297 mod.Data_Mem.F_M.MRAM\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5212_ mod.Data_Mem.F_M.MRAM\[7\]\[4\] mod.Data_Mem.F_M.MRAM\[6\]\[4\] _1876_ _1877_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _1752_ _1748_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5143_ _1651_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7801__I mod.Data_Mem.F_M.MRAM\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5074_ mod.Data_Mem.F_M.MRAM\[3\]\[2\] mod.Data_Mem.F_M.MRAM\[2\]\[2\] _1519_ _1741_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4025_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6417__I _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__I0 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__A2 mod.Data_Mem.F_M.MRAM\[773\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ _2540_ mod.Data_Mem.F_M.MRAM\[789\]\[5\] _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7715_ _3851_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4927_ _1518_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5792__A1 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7646_ mod.Data_Mem.F_M.MRAM\[788\]\[7\] _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4858_ _1521_ _1492_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5544__A1 _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7577_ _3776_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5544__B2 _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4789_ _1330_ _1345_ _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6528_ _2618_ _3129_ _3131_ _2073_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _2722_ mod.Data_Mem.F_M.MRAM\[0\]\[2\] _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5940__B _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8129_ mod.Data_Mem.F_M.out_data\[39\] net40 net275 mod.Arithmetic.CN.I_in\[39\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_87_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4048__S _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6272__A2 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5231__I _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4283__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__A2 mod.Data_Mem.F_M.MRAM\[789\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5387__B _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6062__I _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6011__B _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5406__I _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4310__I _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5838__A2 _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4510__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout180_I net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout278_I net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5141__I _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__A2 mod.Data_Mem.F_M.MRAM\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ _2081_ _2439_ _2453_ _1499_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4026__A1 mod.Arithmetic.CN.I_in\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5074__I0 mod.Data_Mem.F_M.MRAM\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ _2375_ _2377_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7068__I mod.Data_Mem.F_M.MRAM\[20\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7500_ _3728_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4712_ _1365_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8480_ _0576_ net289 mod.Data_Mem.F_M.MRAM\[798\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5692_ _1768_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7431_ mod.Data_Mem.F_M.MRAM\[777\]\[0\] _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5377__I1 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _1063_ _1178_ mod.Arithmetic.CN.I_in\[30\] _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _3654_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4574_ _1125_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _2923_ _2924_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7293_ _3612_ _3606_ _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8469__CLK net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6487__C1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout93_I net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6244_ _2617_ _2857_ _2195_ _2203_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4501__A2 mod.Arithmetic.CN.I_in\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ _2772_ _2789_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ mod.Data_Mem.F_M.MRAM\[786\]\[2\] _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5057_ _1680_ _1723_ _1724_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4008_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__4804__A3 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6006__A2 mod.Data_Mem.F_M.MRAM\[21\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7054__I1 mod.Data_Mem.F_M.MRAM\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4017__A1 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4017__B2 mod.Arithmetic.I_out\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ _2269_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7629_ _2009_ _3804_ _3808_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5368__I1 mod.Data_Mem.F_M.MRAM\[16\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6493__A2 mod.Data_Mem.F_M.MRAM\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5162__S _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_403 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_414 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_425 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_436 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_447 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_458 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_75_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_469 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4256__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7986__CLK net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7985__RN net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5851__S1 _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5359__I1 mod.Data_Mem.F_M.MRAM\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5337__S _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6181__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__I0 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4040__I mod.Arithmetic.I_out\[73\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ _0962_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5287__A3 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4975__I _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8162__RN net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4495__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6236__A2 _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7980_ _0206_ net86 mod.Data_Mem.F_M.MRAM\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5295__I0 mod.Data_Mem.F_M.MRAM\[771\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6931_ _3242_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4798__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5995__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4924__B _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7036__I1 mod.Data_Mem.F_M.MRAM\[18\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _3353_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5813_ _2426_ _2429_ _2430_ _2431_ _2436_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6793_ net7 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8532_ _0036_ net252 mod.Data_Mem.F_M.out_data\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5744_ _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8463_ _0559_ net321 mod.Data_Mem.F_M.MRAM\[795\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5675_ _2304_ mod.Data_Mem.F_M.MRAM\[796\]\[3\] _2254_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7414_ _3680_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _1293_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8394_ _0490_ net201 mod.Data_Mem.F_M.MRAM\[786\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7345_ _3645_ mod.Data_Mem.F_M.MRAM\[771\]\[5\] _3643_ _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4557_ _0633_ mod.Arithmetic.CN.I_in\[53\] _1114_ _1116_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7276_ _3600_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4488_ _1048_ _1077_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4885__I _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _2165_ _1836_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _1607_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6227__A2 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _1769_ _1775_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4238__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6089_ _2705_ mod.Data_Mem.F_M.MRAM\[790\]\[0\] mod.Data_Mem.F_M.MRAM\[791\]\[0\]
+ _2115_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5986__A1 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__A1 _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3964__I _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6163__A1 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5210__I0 mod.Data_Mem.F_M.MRAM\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5910__A1 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 net6 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__A1 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__A2 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8164__CLK net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7018__I1 mod.Data_Mem.F_M.MRAM\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout143_I net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5067__S _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout310_I net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5460_ _2106_ _2108_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _0988_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4704__A2 mod.Arithmetic.ACTI.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5901__A1 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _2052_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5752__I1 mod.Data_Mem.F_M.MRAM\[783\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7130_ _3450_ mod.Data_Mem.F_M.MRAM\[19\]\[1\] _3513_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4342_ _1007_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout308 net309 net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__6457__A2 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout319 net324 net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__8135__RN net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7061_ _3477_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6701__I0 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4273_ _0868_ _0888_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6012_ _2183_ _2146_ _2630_ _2258_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

