VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tiny_user_project
  CLASS BLOCK ;
  FOREIGN tiny_user_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 700.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 483.840 4.000 484.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 490.560 4.000 491.120 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 241.920 4.000 242.480 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 423.360 4.000 423.920 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.960 4.000 289.520 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.640 4.000 249.200 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 696.000 370.160 699.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 141.120 699.000 141.680 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 658.560 699.000 659.120 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 696.000 470.960 699.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 1.000 686.000 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 696.000 87.920 699.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 696.000 558.320 699.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 1.000 491.120 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 698.880 696.000 699.440 699.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 604.800 699.000 605.360 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 1.000 578.480 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 1.000 94.640 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 584.640 4.000 585.200 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 477.120 4.000 477.680 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 544.320 4.000 544.880 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 436.800 4.000 437.360 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 692.160 699.000 692.720 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 1.000 457.520 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 295.680 4.000 296.240 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 1.000 591.920 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 73.920 4.000 74.480 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 624.960 4.000 625.520 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 696.000 625.520 699.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 618.240 699.000 618.800 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 530.880 699.000 531.440 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 685.440 699.000 686.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 315.840 699.000 316.400 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 134.400 4.000 134.960 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 134.400 699.000 134.960 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 696.000 571.760 699.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 322.560 4.000 323.120 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 362.880 4.000 363.440 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 490.560 699.000 491.120 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 450.240 699.000 450.800 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 696.000 27.440 699.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 1.000 430.640 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 181.440 4.000 182.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 1.000 638.960 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 696.000 444.080 699.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 1.000 202.160 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 1.000 67.760 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 696.000 34.160 699.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 696.000 249.200 699.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 696.000 188.720 699.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 696.000 403.760 699.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 1.000 598.640 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 181.440 699.000 182.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 696.000 679.280 699.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 201.600 4.000 202.160 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 100.800 4.000 101.360 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 638.400 4.000 638.960 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 1.000 585.200 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 696.000 14.000 699.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 356.160 699.000 356.720 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 268.800 699.000 269.360 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 1.000 659.120 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 215.040 4.000 215.600 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 696.000 612.080 699.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 114.240 699.000 114.800 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 571.200 4.000 571.760 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 631.680 699.000 632.240 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 696.000 390.320 699.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 282.240 699.000 282.800 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 524.160 4.000 524.720 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 94.080 4.000 94.640 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 696.000 511.280 699.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 551.040 4.000 551.600 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 696.000 336.560 699.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 349.440 4.000 350.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 678.720 699.000 679.280 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 696.000 114.800 699.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 696.000 215.600 699.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 1.000 450.800 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 696.000 686.000 699.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 698.880 4.000 699.440 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 517.440 4.000 518.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 1.000 282.800 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 584.640 699.000 585.200 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 1.000 81.200 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 1.000 652.400 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 696.000 155.120 699.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 1.000 47.600 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 67.200 699.000 67.760 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 463.680 4.000 464.240 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 154.560 699.000 155.120 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 262.080 4.000 262.640 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 1.000 612.080 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 20.160 699.000 20.720 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 1.000 296.240 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 1.000 235.760 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 696.000 491.120 699.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 1.000 477.680 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 248.640 699.000 249.200 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 696.000 638.960 699.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 1.000 249.200 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 696.000 437.360 699.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 255.360 4.000 255.920 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 1.000 464.240 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 1.000 417.200 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 1.000 168.560 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 33.600 4.000 34.160 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 696.000 323.120 699.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 322.560 1.000 323.120 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 696.000 296.240 699.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 127.680 4.000 128.240 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 396.480 4.000 397.040 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 1.000 511.280 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 1.000 182.000 4.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 356.160 4.000 356.720 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 651.840 699.000 652.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 309.120 699.000 309.680 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 1.000 215.600 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 696.000 282.800 699.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 611.520 4.000 612.080 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 504.000 699.000 504.560 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 696.000 67.760 699.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 107.520 699.000 108.080 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 696.000 350.000 699.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 107.520 4.000 108.080 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 696.000 161.840 699.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 147.840 699.000 148.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 530.880 4.000 531.440 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 309.120 4.000 309.680 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 524.160 699.000 524.720 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 696.000 356.720 699.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 696.000 148.400 699.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 696.000 430.640 699.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 631.680 4.000 632.240 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 658.560 4.000 659.120 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 174.720 699.000 175.280 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 696.000 309.680 699.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 53.760 4.000 54.320 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 696.000 591.920 699.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 282.240 4.000 282.800 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 470.400 4.000 470.960 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 696.000 54.320 699.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 618.240 4.000 618.800 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 1.000 497.840 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 685.440 4.000 686.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 1.000 316.400 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 696.000 383.600 699.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 383.040 699.000 383.600 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 1.000 242.480 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 1.000 336.560 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 235.200 4.000 235.760 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 696.000 659.120 699.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 6.720 699.000 7.280 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 1.000 229.040 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 510.720 699.000 511.280 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 1.000 437.360 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 696.000 329.840 699.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 696.000 269.360 699.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 696.000 61.040 699.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 696.000 276.080 699.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 1.000 329.840 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 235.200 699.000 235.760 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 696.000 544.880 699.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.280 696.000 497.840 699.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 188.160 4.000 188.720 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 208.320 4.000 208.880 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 696.000 20.720 699.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 1.000 255.920 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 638.400 699.000 638.960 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 1.000 121.520 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 463.680 699.000 464.240 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 20.160 4.000 20.720 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 1.000 410.480 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 696.000 182.000 699.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 1.000 141.680 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 255.360 699.000 255.920 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 13.440 4.000 14.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 696.000 632.240 699.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 696.000 605.360 699.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 376.320 699.000 376.880 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.880 4.000 27.440 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 504.000 4.000 504.560 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 1.000 262.640 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 288.960 699.000 289.520 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 598.080 4.000 598.640 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 389.760 699.000 390.320 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 696.000 343.280 699.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 577.920 699.000 578.480 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 1.000 370.160 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 329.280 699.000 329.840 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 100.800 699.000 101.360 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 692.160 4.000 692.720 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 436.800 699.000 437.360 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 1.000 208.880 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 315.840 4.000 316.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 1.000 376.880 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 678.720 4.000 679.280 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 696.000 423.920 699.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 557.760 699.000 558.320 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 1.000 302.960 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 161.280 4.000 161.840 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 322.560 699.000 323.120 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 33.600 699.000 34.160 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 696.000 410.480 699.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 127.680 699.000 128.240 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 1.000 343.280 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 696.000 376.880 699.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 564.480 699.000 565.040 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 275.520 699.000 276.080 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 13.440 699.000 14.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 94.080 699.000 94.640 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 114.240 4.000 114.800 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 1.000 679.280 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 215.040 699.000 215.600 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 591.360 699.000 591.920 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 1.000 40.880 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 1.000 289.520 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 696.000 108.080 699.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 696.000 101.360 699.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 497.280 4.000 497.840 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 1.000 161.840 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 631.680 1.000 632.240 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 696.000 397.040 699.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 696.000 242.480 699.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 672.000 4.000 672.560 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 47.040 699.000 47.600 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 665.280 4.000 665.840 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 477.120 699.000 477.680 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 696.000 262.640 699.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 168.000 699.000 168.560 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 696.000 531.440 699.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 483.840 699.000 484.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 268.800 4.000 269.360 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 416.640 699.000 417.200 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 696.000 565.040 699.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 1.000 188.720 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 1.000 605.360 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 53.760 699.000 54.320 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 201.600 699.000 202.160 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 696.000 672.560 699.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 40.320 4.000 40.880 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 336.000 699.000 336.560 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 262.080 699.000 262.640 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 497.280 699.000 497.840 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 396.480 699.000 397.040 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 696.000 7.280 699.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 557.760 4.000 558.320 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 1.000 518.000 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 1.000 618.800 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 1.000 101.360 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 87.360 4.000 87.920 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 696.000 47.600 699.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 60.480 699.000 61.040 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 696.000 134.960 699.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 409.920 4.000 410.480 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 696.000 289.520 699.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 696.000 518.000 699.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 1.000 195.440 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 430.080 699.000 430.640 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 1.000 625.520 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 696.000 141.680 699.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 1.000 128.240 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 430.080 4.000 430.640 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 665.280 699.000 665.840 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 696.000 692.720 699.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 598.080 699.000 598.640 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 696.000 302.960 699.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 571.200 699.000 571.760 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 1.000 356.720 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 696.000 121.520 699.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 1.000 20.720 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 1.000 7.280 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 696.000 94.640 699.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 1.000 363.440 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 302.400 4.000 302.960 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 383.040 4.000 383.600 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 87.360 699.000 87.920 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 696.000 255.920 699.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 443.520 4.000 444.080 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 1.000 134.960 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 1.000 309.680 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 696.000 578.480 699.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 1.000 558.320 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 80.640 4.000 81.200 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 510.720 4.000 511.280 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 6.720 4.000 7.280 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 651.840 4.000 652.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 1.000 538.160 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 696.000 229.040 699.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 1.000 692.720 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 443.520 699.000 444.080 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 376.320 4.000 376.880 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 362.880 699.000 363.440 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 1.000 531.440 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 696.000 618.800 699.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 73.920 699.000 74.480 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 696.000 417.200 699.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 1.000 645.680 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 342.720 4.000 343.280 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 1.000 87.920 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 349.440 699.000 350.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 168.000 4.000 168.560 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 456.960 699.000 457.520 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 1.000 175.280 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 1.000 665.840 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 696.000 202.160 699.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 696.000 598.640 699.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 537.600 699.000 538.160 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 696.000 175.280 699.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 450.240 4.000 450.800 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 682.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 682.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 120.960 699.000 121.520 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 696.000 128.240 699.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 241.920 699.000 242.480 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 696.000 464.240 699.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 696.000 316.400 699.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 403.200 4.000 403.760 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 1.000 61.040 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 389.760 1.000 390.320 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 67.200 4.000 67.760 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 470.400 699.000 470.960 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 1.000 444.080 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 389.760 4.000 390.320 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 221.760 699.000 222.320 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.000 1.000 672.560 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 47.040 4.000 47.600 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 696.000 652.400 699.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 1.000 397.040 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 564.480 1.000 565.040 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 161.280 699.000 161.840 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 696.000 81.200 699.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 120.960 4.000 121.520 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 1.000 74.480 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 696.000 235.760 699.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 409.920 699.000 410.480 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 672.000 699.000 672.560 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 1.000 276.080 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 275.520 4.000 276.080 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 295.680 699.000 296.240 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 1.000 544.880 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 696.000 538.160 699.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 1.000 524.720 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 174.720 4.000 175.280 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 1.000 34.160 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 0.000 699.000 0.560 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 188.160 699.000 188.720 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 696.000 222.320 699.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 611.520 699.000 612.080 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 537.600 4.000 538.160 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 591.360 4.000 591.920 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 564.480 4.000 565.040 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 1.000 27.440 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 147.840 4.000 148.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 369.600 699.000 370.160 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 1.000 403.760 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 696.000 477.680 699.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 696.000 645.680 699.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 696.000 40.880 699.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 1.000 108.080 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 329.280 4.000 329.840 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 696.000 665.840 699.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 416.640 4.000 417.200 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 551.040 699.000 551.600 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 228.480 699.000 229.040 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 1.000 484.400 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 696.000 585.200 699.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 696.000 168.560 699.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1.000 222.320 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 423.360 699.000 423.920 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 1.000 571.760 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 208.320 699.000 208.880 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 369.600 4.000 370.160 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 26.880 699.000 27.440 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 1.000 114.800 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 1.000 350.000 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 302.400 699.000 302.960 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 696.000 551.600 699.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 624.960 699.000 625.520 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 40.320 699.000 40.880 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 141.120 4.000 141.680 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 403.200 699.000 403.760 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 1.000 14.000 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 645.120 699.000 645.680 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.160 696.000 524.720 699.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 80.640 699.000 81.200 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 696.000 504.560 699.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 194.880 4.000 195.440 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 221.760 4.000 222.320 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 1.000 470.960 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 1.000 551.600 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 336.000 4.000 336.560 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 604.800 4.000 605.360 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 696.000 195.440 699.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 228.480 4.000 229.040 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 1.000 148.400 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 1.000 54.320 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 362.880 696.000 363.440 699.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 696.000 208.880 699.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 1.000 383.600 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 696.000 484.400 699.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 194.880 699.000 195.440 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 456.960 4.000 457.520 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 544.320 699.000 544.880 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 1.000 155.120 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 1.000 269.360 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 60.480 4.000 61.040 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 517.440 699.000 518.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 1.000 423.920 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 456.960 696.000 457.520 699.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 696.000 450.800 699.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 645.120 4.000 645.680 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 696.000 74.480 699.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 1.000 504.560 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 154.560 4.000 155.120 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 577.920 4.000 578.480 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 696.000 342.720 699.000 343.280 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 693.280 685.290 ;
      LAYER Metal2 ;
        RECT 0.140 699.300 698.180 699.350 ;
        RECT 0.140 695.700 6.420 699.300 ;
        RECT 7.580 695.700 13.140 699.300 ;
        RECT 14.300 695.700 19.860 699.300 ;
        RECT 21.020 695.700 26.580 699.300 ;
        RECT 27.740 695.700 33.300 699.300 ;
        RECT 34.460 695.700 40.020 699.300 ;
        RECT 41.180 695.700 46.740 699.300 ;
        RECT 47.900 695.700 53.460 699.300 ;
        RECT 54.620 695.700 60.180 699.300 ;
        RECT 61.340 695.700 66.900 699.300 ;
        RECT 68.060 695.700 73.620 699.300 ;
        RECT 74.780 695.700 80.340 699.300 ;
        RECT 81.500 695.700 87.060 699.300 ;
        RECT 88.220 695.700 93.780 699.300 ;
        RECT 94.940 695.700 100.500 699.300 ;
        RECT 101.660 695.700 107.220 699.300 ;
        RECT 108.380 695.700 113.940 699.300 ;
        RECT 115.100 695.700 120.660 699.300 ;
        RECT 121.820 695.700 127.380 699.300 ;
        RECT 128.540 695.700 134.100 699.300 ;
        RECT 135.260 695.700 140.820 699.300 ;
        RECT 141.980 695.700 147.540 699.300 ;
        RECT 148.700 695.700 154.260 699.300 ;
        RECT 155.420 695.700 160.980 699.300 ;
        RECT 162.140 695.700 167.700 699.300 ;
        RECT 168.860 695.700 174.420 699.300 ;
        RECT 175.580 695.700 181.140 699.300 ;
        RECT 182.300 695.700 187.860 699.300 ;
        RECT 189.020 695.700 194.580 699.300 ;
        RECT 195.740 695.700 201.300 699.300 ;
        RECT 202.460 695.700 208.020 699.300 ;
        RECT 209.180 695.700 214.740 699.300 ;
        RECT 215.900 695.700 221.460 699.300 ;
        RECT 222.620 695.700 228.180 699.300 ;
        RECT 229.340 695.700 234.900 699.300 ;
        RECT 236.060 695.700 241.620 699.300 ;
        RECT 242.780 695.700 248.340 699.300 ;
        RECT 249.500 695.700 255.060 699.300 ;
        RECT 256.220 695.700 261.780 699.300 ;
        RECT 262.940 695.700 268.500 699.300 ;
        RECT 269.660 695.700 275.220 699.300 ;
        RECT 276.380 695.700 281.940 699.300 ;
        RECT 283.100 695.700 288.660 699.300 ;
        RECT 289.820 695.700 295.380 699.300 ;
        RECT 296.540 695.700 302.100 699.300 ;
        RECT 303.260 695.700 308.820 699.300 ;
        RECT 309.980 695.700 315.540 699.300 ;
        RECT 316.700 695.700 322.260 699.300 ;
        RECT 323.420 695.700 328.980 699.300 ;
        RECT 330.140 695.700 335.700 699.300 ;
        RECT 336.860 695.700 342.420 699.300 ;
        RECT 343.580 695.700 349.140 699.300 ;
        RECT 350.300 695.700 355.860 699.300 ;
        RECT 357.020 695.700 362.580 699.300 ;
        RECT 363.740 695.700 369.300 699.300 ;
        RECT 370.460 695.700 376.020 699.300 ;
        RECT 377.180 695.700 382.740 699.300 ;
        RECT 383.900 695.700 389.460 699.300 ;
        RECT 390.620 695.700 396.180 699.300 ;
        RECT 397.340 695.700 402.900 699.300 ;
        RECT 404.060 695.700 409.620 699.300 ;
        RECT 410.780 695.700 416.340 699.300 ;
        RECT 417.500 695.700 423.060 699.300 ;
        RECT 424.220 695.700 429.780 699.300 ;
        RECT 430.940 695.700 436.500 699.300 ;
        RECT 437.660 695.700 443.220 699.300 ;
        RECT 444.380 695.700 449.940 699.300 ;
        RECT 451.100 695.700 456.660 699.300 ;
        RECT 457.820 695.700 463.380 699.300 ;
        RECT 464.540 695.700 470.100 699.300 ;
        RECT 471.260 695.700 476.820 699.300 ;
        RECT 477.980 695.700 483.540 699.300 ;
        RECT 484.700 695.700 490.260 699.300 ;
        RECT 491.420 695.700 496.980 699.300 ;
        RECT 498.140 695.700 503.700 699.300 ;
        RECT 504.860 695.700 510.420 699.300 ;
        RECT 511.580 695.700 517.140 699.300 ;
        RECT 518.300 695.700 523.860 699.300 ;
        RECT 525.020 695.700 530.580 699.300 ;
        RECT 531.740 695.700 537.300 699.300 ;
        RECT 538.460 695.700 544.020 699.300 ;
        RECT 545.180 695.700 550.740 699.300 ;
        RECT 551.900 695.700 557.460 699.300 ;
        RECT 558.620 695.700 564.180 699.300 ;
        RECT 565.340 695.700 570.900 699.300 ;
        RECT 572.060 695.700 577.620 699.300 ;
        RECT 578.780 695.700 584.340 699.300 ;
        RECT 585.500 695.700 591.060 699.300 ;
        RECT 592.220 695.700 597.780 699.300 ;
        RECT 598.940 695.700 604.500 699.300 ;
        RECT 605.660 695.700 611.220 699.300 ;
        RECT 612.380 695.700 617.940 699.300 ;
        RECT 619.100 695.700 624.660 699.300 ;
        RECT 625.820 695.700 631.380 699.300 ;
        RECT 632.540 695.700 638.100 699.300 ;
        RECT 639.260 695.700 644.820 699.300 ;
        RECT 645.980 695.700 651.540 699.300 ;
        RECT 652.700 695.700 658.260 699.300 ;
        RECT 659.420 695.700 664.980 699.300 ;
        RECT 666.140 695.700 671.700 699.300 ;
        RECT 672.860 695.700 678.420 699.300 ;
        RECT 679.580 695.700 685.140 699.300 ;
        RECT 686.300 695.700 691.860 699.300 ;
        RECT 693.020 695.700 698.180 699.300 ;
        RECT 0.140 4.300 698.180 695.700 ;
        RECT 0.860 4.000 6.420 4.300 ;
        RECT 7.580 4.000 13.140 4.300 ;
        RECT 14.300 4.000 19.860 4.300 ;
        RECT 21.020 4.000 26.580 4.300 ;
        RECT 27.740 4.000 33.300 4.300 ;
        RECT 34.460 4.000 40.020 4.300 ;
        RECT 41.180 4.000 46.740 4.300 ;
        RECT 47.900 4.000 53.460 4.300 ;
        RECT 54.620 4.000 60.180 4.300 ;
        RECT 61.340 4.000 66.900 4.300 ;
        RECT 68.060 4.000 73.620 4.300 ;
        RECT 74.780 4.000 80.340 4.300 ;
        RECT 81.500 4.000 87.060 4.300 ;
        RECT 88.220 4.000 93.780 4.300 ;
        RECT 94.940 4.000 100.500 4.300 ;
        RECT 101.660 4.000 107.220 4.300 ;
        RECT 108.380 4.000 113.940 4.300 ;
        RECT 115.100 4.000 120.660 4.300 ;
        RECT 121.820 4.000 127.380 4.300 ;
        RECT 128.540 4.000 134.100 4.300 ;
        RECT 135.260 4.000 140.820 4.300 ;
        RECT 141.980 4.000 147.540 4.300 ;
        RECT 148.700 4.000 154.260 4.300 ;
        RECT 155.420 4.000 160.980 4.300 ;
        RECT 162.140 4.000 167.700 4.300 ;
        RECT 168.860 4.000 174.420 4.300 ;
        RECT 175.580 4.000 181.140 4.300 ;
        RECT 182.300 4.000 187.860 4.300 ;
        RECT 189.020 4.000 194.580 4.300 ;
        RECT 195.740 4.000 201.300 4.300 ;
        RECT 202.460 4.000 208.020 4.300 ;
        RECT 209.180 4.000 214.740 4.300 ;
        RECT 215.900 4.000 221.460 4.300 ;
        RECT 222.620 4.000 228.180 4.300 ;
        RECT 229.340 4.000 234.900 4.300 ;
        RECT 236.060 4.000 241.620 4.300 ;
        RECT 242.780 4.000 248.340 4.300 ;
        RECT 249.500 4.000 255.060 4.300 ;
        RECT 256.220 4.000 261.780 4.300 ;
        RECT 262.940 4.000 268.500 4.300 ;
        RECT 269.660 4.000 275.220 4.300 ;
        RECT 276.380 4.000 281.940 4.300 ;
        RECT 283.100 4.000 288.660 4.300 ;
        RECT 289.820 4.000 295.380 4.300 ;
        RECT 296.540 4.000 302.100 4.300 ;
        RECT 303.260 4.000 308.820 4.300 ;
        RECT 309.980 4.000 315.540 4.300 ;
        RECT 316.700 4.000 322.260 4.300 ;
        RECT 323.420 4.000 328.980 4.300 ;
        RECT 330.140 4.000 335.700 4.300 ;
        RECT 336.860 4.000 342.420 4.300 ;
        RECT 343.580 4.000 349.140 4.300 ;
        RECT 350.300 4.000 355.860 4.300 ;
        RECT 357.020 4.000 362.580 4.300 ;
        RECT 363.740 4.000 369.300 4.300 ;
        RECT 370.460 4.000 376.020 4.300 ;
        RECT 377.180 4.000 382.740 4.300 ;
        RECT 383.900 4.000 389.460 4.300 ;
        RECT 390.620 4.000 396.180 4.300 ;
        RECT 397.340 4.000 402.900 4.300 ;
        RECT 404.060 4.000 409.620 4.300 ;
        RECT 410.780 4.000 416.340 4.300 ;
        RECT 417.500 4.000 423.060 4.300 ;
        RECT 424.220 4.000 429.780 4.300 ;
        RECT 430.940 4.000 436.500 4.300 ;
        RECT 437.660 4.000 443.220 4.300 ;
        RECT 444.380 4.000 449.940 4.300 ;
        RECT 451.100 4.000 456.660 4.300 ;
        RECT 457.820 4.000 463.380 4.300 ;
        RECT 464.540 4.000 470.100 4.300 ;
        RECT 471.260 4.000 476.820 4.300 ;
        RECT 477.980 4.000 483.540 4.300 ;
        RECT 484.700 4.000 490.260 4.300 ;
        RECT 491.420 4.000 496.980 4.300 ;
        RECT 498.140 4.000 503.700 4.300 ;
        RECT 504.860 4.000 510.420 4.300 ;
        RECT 511.580 4.000 517.140 4.300 ;
        RECT 518.300 4.000 523.860 4.300 ;
        RECT 525.020 4.000 530.580 4.300 ;
        RECT 531.740 4.000 537.300 4.300 ;
        RECT 538.460 4.000 544.020 4.300 ;
        RECT 545.180 4.000 550.740 4.300 ;
        RECT 551.900 4.000 557.460 4.300 ;
        RECT 558.620 4.000 564.180 4.300 ;
        RECT 565.340 4.000 570.900 4.300 ;
        RECT 572.060 4.000 577.620 4.300 ;
        RECT 578.780 4.000 584.340 4.300 ;
        RECT 585.500 4.000 591.060 4.300 ;
        RECT 592.220 4.000 597.780 4.300 ;
        RECT 598.940 4.000 604.500 4.300 ;
        RECT 605.660 4.000 611.220 4.300 ;
        RECT 612.380 4.000 617.940 4.300 ;
        RECT 619.100 4.000 624.660 4.300 ;
        RECT 625.820 4.000 631.380 4.300 ;
        RECT 632.540 4.000 638.100 4.300 ;
        RECT 639.260 4.000 644.820 4.300 ;
        RECT 645.980 4.000 651.540 4.300 ;
        RECT 652.700 4.000 658.260 4.300 ;
        RECT 659.420 4.000 664.980 4.300 ;
        RECT 666.140 4.000 671.700 4.300 ;
        RECT 672.860 4.000 678.420 4.300 ;
        RECT 679.580 4.000 685.140 4.300 ;
        RECT 686.300 4.000 691.860 4.300 ;
        RECT 693.020 4.000 698.180 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 698.580 0.700 699.300 ;
        RECT 4.300 698.580 698.230 699.300 ;
        RECT 0.090 693.020 698.230 698.580 ;
        RECT 0.090 691.860 0.700 693.020 ;
        RECT 4.300 691.860 695.700 693.020 ;
        RECT 0.090 686.300 698.230 691.860 ;
        RECT 0.090 685.140 0.700 686.300 ;
        RECT 4.300 685.140 695.700 686.300 ;
        RECT 0.090 679.580 698.230 685.140 ;
        RECT 0.090 678.420 0.700 679.580 ;
        RECT 4.300 678.420 695.700 679.580 ;
        RECT 0.090 672.860 698.230 678.420 ;
        RECT 0.090 671.700 0.700 672.860 ;
        RECT 4.300 671.700 695.700 672.860 ;
        RECT 0.090 666.140 698.230 671.700 ;
        RECT 0.090 664.980 0.700 666.140 ;
        RECT 4.300 664.980 695.700 666.140 ;
        RECT 0.090 659.420 698.230 664.980 ;
        RECT 0.090 658.260 0.700 659.420 ;
        RECT 4.300 658.260 695.700 659.420 ;
        RECT 0.090 652.700 698.230 658.260 ;
        RECT 0.090 651.540 0.700 652.700 ;
        RECT 4.300 651.540 695.700 652.700 ;
        RECT 0.090 645.980 698.230 651.540 ;
        RECT 0.090 644.820 0.700 645.980 ;
        RECT 4.300 644.820 695.700 645.980 ;
        RECT 0.090 639.260 698.230 644.820 ;
        RECT 0.090 638.100 0.700 639.260 ;
        RECT 4.300 638.100 695.700 639.260 ;
        RECT 0.090 632.540 698.230 638.100 ;
        RECT 0.090 631.380 0.700 632.540 ;
        RECT 4.300 631.380 695.700 632.540 ;
        RECT 0.090 625.820 698.230 631.380 ;
        RECT 0.090 624.660 0.700 625.820 ;
        RECT 4.300 624.660 695.700 625.820 ;
        RECT 0.090 619.100 698.230 624.660 ;
        RECT 0.090 617.940 0.700 619.100 ;
        RECT 4.300 617.940 695.700 619.100 ;
        RECT 0.090 612.380 698.230 617.940 ;
        RECT 0.090 611.220 0.700 612.380 ;
        RECT 4.300 611.220 695.700 612.380 ;
        RECT 0.090 605.660 698.230 611.220 ;
        RECT 0.090 604.500 0.700 605.660 ;
        RECT 4.300 604.500 695.700 605.660 ;
        RECT 0.090 598.940 698.230 604.500 ;
        RECT 0.090 597.780 0.700 598.940 ;
        RECT 4.300 597.780 695.700 598.940 ;
        RECT 0.090 592.220 698.230 597.780 ;
        RECT 0.090 591.060 0.700 592.220 ;
        RECT 4.300 591.060 695.700 592.220 ;
        RECT 0.090 585.500 698.230 591.060 ;
        RECT 0.090 584.340 0.700 585.500 ;
        RECT 4.300 584.340 695.700 585.500 ;
        RECT 0.090 578.780 698.230 584.340 ;
        RECT 0.090 577.620 0.700 578.780 ;
        RECT 4.300 577.620 695.700 578.780 ;
        RECT 0.090 572.060 698.230 577.620 ;
        RECT 0.090 570.900 0.700 572.060 ;
        RECT 4.300 570.900 695.700 572.060 ;
        RECT 0.090 565.340 698.230 570.900 ;
        RECT 0.090 564.180 0.700 565.340 ;
        RECT 4.300 564.180 695.700 565.340 ;
        RECT 0.090 558.620 698.230 564.180 ;
        RECT 0.090 557.460 0.700 558.620 ;
        RECT 4.300 557.460 695.700 558.620 ;
        RECT 0.090 551.900 698.230 557.460 ;
        RECT 0.090 550.740 0.700 551.900 ;
        RECT 4.300 550.740 695.700 551.900 ;
        RECT 0.090 545.180 698.230 550.740 ;
        RECT 0.090 544.020 0.700 545.180 ;
        RECT 4.300 544.020 695.700 545.180 ;
        RECT 0.090 538.460 698.230 544.020 ;
        RECT 0.090 537.300 0.700 538.460 ;
        RECT 4.300 537.300 695.700 538.460 ;
        RECT 0.090 531.740 698.230 537.300 ;
        RECT 0.090 530.580 0.700 531.740 ;
        RECT 4.300 530.580 695.700 531.740 ;
        RECT 0.090 525.020 698.230 530.580 ;
        RECT 0.090 523.860 0.700 525.020 ;
        RECT 4.300 523.860 695.700 525.020 ;
        RECT 0.090 518.300 698.230 523.860 ;
        RECT 0.090 517.140 0.700 518.300 ;
        RECT 4.300 517.140 695.700 518.300 ;
        RECT 0.090 511.580 698.230 517.140 ;
        RECT 0.090 510.420 0.700 511.580 ;
        RECT 4.300 510.420 695.700 511.580 ;
        RECT 0.090 504.860 698.230 510.420 ;
        RECT 0.090 503.700 0.700 504.860 ;
        RECT 4.300 503.700 695.700 504.860 ;
        RECT 0.090 498.140 698.230 503.700 ;
        RECT 0.090 496.980 0.700 498.140 ;
        RECT 4.300 496.980 695.700 498.140 ;
        RECT 0.090 491.420 698.230 496.980 ;
        RECT 0.090 490.260 0.700 491.420 ;
        RECT 4.300 490.260 695.700 491.420 ;
        RECT 0.090 484.700 698.230 490.260 ;
        RECT 0.090 483.540 0.700 484.700 ;
        RECT 4.300 483.540 695.700 484.700 ;
        RECT 0.090 477.980 698.230 483.540 ;
        RECT 0.090 476.820 0.700 477.980 ;
        RECT 4.300 476.820 695.700 477.980 ;
        RECT 0.090 471.260 698.230 476.820 ;
        RECT 0.090 470.100 0.700 471.260 ;
        RECT 4.300 470.100 695.700 471.260 ;
        RECT 0.090 464.540 698.230 470.100 ;
        RECT 0.090 463.380 0.700 464.540 ;
        RECT 4.300 463.380 695.700 464.540 ;
        RECT 0.090 457.820 698.230 463.380 ;
        RECT 0.090 456.660 0.700 457.820 ;
        RECT 4.300 456.660 695.700 457.820 ;
        RECT 0.090 451.100 698.230 456.660 ;
        RECT 0.090 449.940 0.700 451.100 ;
        RECT 4.300 449.940 695.700 451.100 ;
        RECT 0.090 444.380 698.230 449.940 ;
        RECT 0.090 443.220 0.700 444.380 ;
        RECT 4.300 443.220 695.700 444.380 ;
        RECT 0.090 437.660 698.230 443.220 ;
        RECT 0.090 436.500 0.700 437.660 ;
        RECT 4.300 436.500 695.700 437.660 ;
        RECT 0.090 430.940 698.230 436.500 ;
        RECT 0.090 429.780 0.700 430.940 ;
        RECT 4.300 429.780 695.700 430.940 ;
        RECT 0.090 424.220 698.230 429.780 ;
        RECT 0.090 423.060 0.700 424.220 ;
        RECT 4.300 423.060 695.700 424.220 ;
        RECT 0.090 417.500 698.230 423.060 ;
        RECT 0.090 416.340 0.700 417.500 ;
        RECT 4.300 416.340 695.700 417.500 ;
        RECT 0.090 410.780 698.230 416.340 ;
        RECT 0.090 409.620 0.700 410.780 ;
        RECT 4.300 409.620 695.700 410.780 ;
        RECT 0.090 404.060 698.230 409.620 ;
        RECT 0.090 402.900 0.700 404.060 ;
        RECT 4.300 402.900 695.700 404.060 ;
        RECT 0.090 397.340 698.230 402.900 ;
        RECT 0.090 396.180 0.700 397.340 ;
        RECT 4.300 396.180 695.700 397.340 ;
        RECT 0.090 390.620 698.230 396.180 ;
        RECT 0.090 389.460 0.700 390.620 ;
        RECT 4.300 389.460 695.700 390.620 ;
        RECT 0.090 383.900 698.230 389.460 ;
        RECT 0.090 382.740 0.700 383.900 ;
        RECT 4.300 382.740 695.700 383.900 ;
        RECT 0.090 377.180 698.230 382.740 ;
        RECT 0.090 376.020 0.700 377.180 ;
        RECT 4.300 376.020 695.700 377.180 ;
        RECT 0.090 370.460 698.230 376.020 ;
        RECT 0.090 369.300 0.700 370.460 ;
        RECT 4.300 369.300 695.700 370.460 ;
        RECT 0.090 363.740 698.230 369.300 ;
        RECT 0.090 362.580 0.700 363.740 ;
        RECT 4.300 362.580 695.700 363.740 ;
        RECT 0.090 357.020 698.230 362.580 ;
        RECT 0.090 355.860 0.700 357.020 ;
        RECT 4.300 355.860 695.700 357.020 ;
        RECT 0.090 350.300 698.230 355.860 ;
        RECT 0.090 349.140 0.700 350.300 ;
        RECT 4.300 349.140 695.700 350.300 ;
        RECT 0.090 343.580 698.230 349.140 ;
        RECT 0.090 342.420 0.700 343.580 ;
        RECT 4.300 342.420 695.700 343.580 ;
        RECT 0.090 336.860 698.230 342.420 ;
        RECT 0.090 335.700 0.700 336.860 ;
        RECT 4.300 335.700 695.700 336.860 ;
        RECT 0.090 330.140 698.230 335.700 ;
        RECT 0.090 328.980 0.700 330.140 ;
        RECT 4.300 328.980 695.700 330.140 ;
        RECT 0.090 323.420 698.230 328.980 ;
        RECT 0.090 322.260 0.700 323.420 ;
        RECT 4.300 322.260 695.700 323.420 ;
        RECT 0.090 316.700 698.230 322.260 ;
        RECT 0.090 315.540 0.700 316.700 ;
        RECT 4.300 315.540 695.700 316.700 ;
        RECT 0.090 309.980 698.230 315.540 ;
        RECT 0.090 308.820 0.700 309.980 ;
        RECT 4.300 308.820 695.700 309.980 ;
        RECT 0.090 303.260 698.230 308.820 ;
        RECT 0.090 302.100 0.700 303.260 ;
        RECT 4.300 302.100 695.700 303.260 ;
        RECT 0.090 296.540 698.230 302.100 ;
        RECT 0.090 295.380 0.700 296.540 ;
        RECT 4.300 295.380 695.700 296.540 ;
        RECT 0.090 289.820 698.230 295.380 ;
        RECT 0.090 288.660 0.700 289.820 ;
        RECT 4.300 288.660 695.700 289.820 ;
        RECT 0.090 283.100 698.230 288.660 ;
        RECT 0.090 281.940 0.700 283.100 ;
        RECT 4.300 281.940 695.700 283.100 ;
        RECT 0.090 276.380 698.230 281.940 ;
        RECT 0.090 275.220 0.700 276.380 ;
        RECT 4.300 275.220 695.700 276.380 ;
        RECT 0.090 269.660 698.230 275.220 ;
        RECT 0.090 268.500 0.700 269.660 ;
        RECT 4.300 268.500 695.700 269.660 ;
        RECT 0.090 262.940 698.230 268.500 ;
        RECT 0.090 261.780 0.700 262.940 ;
        RECT 4.300 261.780 695.700 262.940 ;
        RECT 0.090 256.220 698.230 261.780 ;
        RECT 0.090 255.060 0.700 256.220 ;
        RECT 4.300 255.060 695.700 256.220 ;
        RECT 0.090 249.500 698.230 255.060 ;
        RECT 0.090 248.340 0.700 249.500 ;
        RECT 4.300 248.340 695.700 249.500 ;
        RECT 0.090 242.780 698.230 248.340 ;
        RECT 0.090 241.620 0.700 242.780 ;
        RECT 4.300 241.620 695.700 242.780 ;
        RECT 0.090 236.060 698.230 241.620 ;
        RECT 0.090 234.900 0.700 236.060 ;
        RECT 4.300 234.900 695.700 236.060 ;
        RECT 0.090 229.340 698.230 234.900 ;
        RECT 0.090 228.180 0.700 229.340 ;
        RECT 4.300 228.180 695.700 229.340 ;
        RECT 0.090 222.620 698.230 228.180 ;
        RECT 0.090 221.460 0.700 222.620 ;
        RECT 4.300 221.460 695.700 222.620 ;
        RECT 0.090 215.900 698.230 221.460 ;
        RECT 0.090 214.740 0.700 215.900 ;
        RECT 4.300 214.740 695.700 215.900 ;
        RECT 0.090 209.180 698.230 214.740 ;
        RECT 0.090 208.020 0.700 209.180 ;
        RECT 4.300 208.020 695.700 209.180 ;
        RECT 0.090 202.460 698.230 208.020 ;
        RECT 0.090 201.300 0.700 202.460 ;
        RECT 4.300 201.300 695.700 202.460 ;
        RECT 0.090 195.740 698.230 201.300 ;
        RECT 0.090 194.580 0.700 195.740 ;
        RECT 4.300 194.580 695.700 195.740 ;
        RECT 0.090 189.020 698.230 194.580 ;
        RECT 0.090 187.860 0.700 189.020 ;
        RECT 4.300 187.860 695.700 189.020 ;
        RECT 0.090 182.300 698.230 187.860 ;
        RECT 0.090 181.140 0.700 182.300 ;
        RECT 4.300 181.140 695.700 182.300 ;
        RECT 0.090 175.580 698.230 181.140 ;
        RECT 0.090 174.420 0.700 175.580 ;
        RECT 4.300 174.420 695.700 175.580 ;
        RECT 0.090 168.860 698.230 174.420 ;
        RECT 0.090 167.700 0.700 168.860 ;
        RECT 4.300 167.700 695.700 168.860 ;
        RECT 0.090 162.140 698.230 167.700 ;
        RECT 0.090 160.980 0.700 162.140 ;
        RECT 4.300 160.980 695.700 162.140 ;
        RECT 0.090 155.420 698.230 160.980 ;
        RECT 0.090 154.260 0.700 155.420 ;
        RECT 4.300 154.260 695.700 155.420 ;
        RECT 0.090 148.700 698.230 154.260 ;
        RECT 0.090 147.540 0.700 148.700 ;
        RECT 4.300 147.540 695.700 148.700 ;
        RECT 0.090 141.980 698.230 147.540 ;
        RECT 0.090 140.820 0.700 141.980 ;
        RECT 4.300 140.820 695.700 141.980 ;
        RECT 0.090 135.260 698.230 140.820 ;
        RECT 0.090 134.100 0.700 135.260 ;
        RECT 4.300 134.100 695.700 135.260 ;
        RECT 0.090 128.540 698.230 134.100 ;
        RECT 0.090 127.380 0.700 128.540 ;
        RECT 4.300 127.380 695.700 128.540 ;
        RECT 0.090 121.820 698.230 127.380 ;
        RECT 0.090 120.660 0.700 121.820 ;
        RECT 4.300 120.660 695.700 121.820 ;
        RECT 0.090 115.100 698.230 120.660 ;
        RECT 0.090 113.940 0.700 115.100 ;
        RECT 4.300 113.940 695.700 115.100 ;
        RECT 0.090 108.380 698.230 113.940 ;
        RECT 0.090 107.220 0.700 108.380 ;
        RECT 4.300 107.220 695.700 108.380 ;
        RECT 0.090 101.660 698.230 107.220 ;
        RECT 0.090 100.500 0.700 101.660 ;
        RECT 4.300 100.500 695.700 101.660 ;
        RECT 0.090 94.940 698.230 100.500 ;
        RECT 0.090 93.780 0.700 94.940 ;
        RECT 4.300 93.780 695.700 94.940 ;
        RECT 0.090 88.220 698.230 93.780 ;
        RECT 0.090 87.060 0.700 88.220 ;
        RECT 4.300 87.060 695.700 88.220 ;
        RECT 0.090 81.500 698.230 87.060 ;
        RECT 0.090 80.340 0.700 81.500 ;
        RECT 4.300 80.340 695.700 81.500 ;
        RECT 0.090 74.780 698.230 80.340 ;
        RECT 0.090 73.620 0.700 74.780 ;
        RECT 4.300 73.620 695.700 74.780 ;
        RECT 0.090 68.060 698.230 73.620 ;
        RECT 0.090 66.900 0.700 68.060 ;
        RECT 4.300 66.900 695.700 68.060 ;
        RECT 0.090 61.340 698.230 66.900 ;
        RECT 0.090 60.180 0.700 61.340 ;
        RECT 4.300 60.180 695.700 61.340 ;
        RECT 0.090 54.620 698.230 60.180 ;
        RECT 0.090 53.460 0.700 54.620 ;
        RECT 4.300 53.460 695.700 54.620 ;
        RECT 0.090 47.900 698.230 53.460 ;
        RECT 0.090 46.740 0.700 47.900 ;
        RECT 4.300 46.740 695.700 47.900 ;
        RECT 0.090 41.180 698.230 46.740 ;
        RECT 0.090 40.020 0.700 41.180 ;
        RECT 4.300 40.020 695.700 41.180 ;
        RECT 0.090 34.460 698.230 40.020 ;
        RECT 0.090 33.300 0.700 34.460 ;
        RECT 4.300 33.300 695.700 34.460 ;
        RECT 0.090 27.740 698.230 33.300 ;
        RECT 0.090 26.580 0.700 27.740 ;
        RECT 4.300 26.580 695.700 27.740 ;
        RECT 0.090 21.020 698.230 26.580 ;
        RECT 0.090 19.860 0.700 21.020 ;
        RECT 4.300 19.860 695.700 21.020 ;
        RECT 0.090 14.300 698.230 19.860 ;
        RECT 0.090 13.140 0.700 14.300 ;
        RECT 4.300 13.140 695.700 14.300 ;
        RECT 0.090 7.580 698.230 13.140 ;
        RECT 0.090 6.420 0.700 7.580 ;
        RECT 4.300 6.420 695.700 7.580 ;
        RECT 0.090 5.180 698.230 6.420 ;
      LAYER Metal4 ;
        RECT 109.900 15.080 175.540 598.550 ;
        RECT 177.740 15.080 252.340 598.550 ;
        RECT 254.540 15.080 329.140 598.550 ;
        RECT 331.340 15.080 405.940 598.550 ;
        RECT 408.140 15.080 482.740 598.550 ;
        RECT 484.940 15.080 559.540 598.550 ;
        RECT 561.740 15.080 636.340 598.550 ;
        RECT 638.540 15.080 692.020 598.550 ;
        RECT 109.900 5.130 692.020 15.080 ;
  END
END tiny_user_project
END LIBRARY

