// This is the unpowered netlist.
module tiny_user_project (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire net574;
 wire net573;
 wire net572;
 wire net571;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire net570;
 wire net569;
 wire net568;
 wire net567;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire net566;
 wire net565;
 wire net564;
 wire net563;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire net395;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net396;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net397;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net433;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net434;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net435;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net463;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net464;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net465;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net466;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net467;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net468;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire \mod.Arithmetic.ACTI.x[0] ;
 wire \mod.Arithmetic.ACTI.x[1] ;
 wire \mod.Arithmetic.ACTI.x[2] ;
 wire \mod.Arithmetic.ACTI.x[3] ;
 wire \mod.Arithmetic.ACTI.x[4] ;
 wire \mod.Arithmetic.ACTI.x[5] ;
 wire \mod.Arithmetic.ACTI.x[6] ;
 wire \mod.Arithmetic.ACTI.x[7] ;
 wire \mod.Arithmetic.CN.F_in[0] ;
 wire \mod.Arithmetic.CN.I_in[10] ;
 wire \mod.Arithmetic.CN.I_in[11] ;
 wire \mod.Arithmetic.CN.I_in[12] ;
 wire \mod.Arithmetic.CN.I_in[13] ;
 wire \mod.Arithmetic.CN.I_in[14] ;
 wire \mod.Arithmetic.CN.I_in[15] ;
 wire \mod.Arithmetic.CN.I_in[16] ;
 wire \mod.Arithmetic.CN.I_in[17] ;
 wire \mod.Arithmetic.CN.I_in[18] ;
 wire \mod.Arithmetic.CN.I_in[19] ;
 wire \mod.Arithmetic.CN.I_in[20] ;
 wire \mod.Arithmetic.CN.I_in[21] ;
 wire \mod.Arithmetic.CN.I_in[22] ;
 wire \mod.Arithmetic.CN.I_in[23] ;
 wire \mod.Arithmetic.CN.I_in[24] ;
 wire \mod.Arithmetic.CN.I_in[25] ;
 wire \mod.Arithmetic.CN.I_in[26] ;
 wire \mod.Arithmetic.CN.I_in[27] ;
 wire \mod.Arithmetic.CN.I_in[28] ;
 wire \mod.Arithmetic.CN.I_in[29] ;
 wire \mod.Arithmetic.CN.I_in[30] ;
 wire \mod.Arithmetic.CN.I_in[31] ;
 wire \mod.Arithmetic.CN.I_in[32] ;
 wire \mod.Arithmetic.CN.I_in[33] ;
 wire \mod.Arithmetic.CN.I_in[34] ;
 wire \mod.Arithmetic.CN.I_in[35] ;
 wire \mod.Arithmetic.CN.I_in[36] ;
 wire \mod.Arithmetic.CN.I_in[37] ;
 wire \mod.Arithmetic.CN.I_in[38] ;
 wire \mod.Arithmetic.CN.I_in[39] ;
 wire \mod.Arithmetic.CN.I_in[40] ;
 wire \mod.Arithmetic.CN.I_in[41] ;
 wire \mod.Arithmetic.CN.I_in[42] ;
 wire \mod.Arithmetic.CN.I_in[43] ;
 wire \mod.Arithmetic.CN.I_in[44] ;
 wire \mod.Arithmetic.CN.I_in[45] ;
 wire \mod.Arithmetic.CN.I_in[46] ;
 wire \mod.Arithmetic.CN.I_in[47] ;
 wire \mod.Arithmetic.CN.I_in[48] ;
 wire \mod.Arithmetic.CN.I_in[49] ;
 wire \mod.Arithmetic.CN.I_in[50] ;
 wire \mod.Arithmetic.CN.I_in[51] ;
 wire \mod.Arithmetic.CN.I_in[52] ;
 wire \mod.Arithmetic.CN.I_in[53] ;
 wire \mod.Arithmetic.CN.I_in[54] ;
 wire \mod.Arithmetic.CN.I_in[55] ;
 wire \mod.Arithmetic.CN.I_in[56] ;
 wire \mod.Arithmetic.CN.I_in[57] ;
 wire \mod.Arithmetic.CN.I_in[58] ;
 wire \mod.Arithmetic.CN.I_in[59] ;
 wire \mod.Arithmetic.CN.I_in[60] ;
 wire \mod.Arithmetic.CN.I_in[61] ;
 wire \mod.Arithmetic.CN.I_in[62] ;
 wire \mod.Arithmetic.CN.I_in[63] ;
 wire \mod.Arithmetic.CN.I_in[64] ;
 wire \mod.Arithmetic.CN.I_in[65] ;
 wire \mod.Arithmetic.CN.I_in[66] ;
 wire \mod.Arithmetic.CN.I_in[67] ;
 wire \mod.Arithmetic.CN.I_in[68] ;
 wire \mod.Arithmetic.CN.I_in[69] ;
 wire \mod.Arithmetic.CN.I_in[70] ;
 wire \mod.Arithmetic.CN.I_in[71] ;
 wire \mod.Arithmetic.CN.I_in[8] ;
 wire \mod.Arithmetic.CN.I_in[9] ;
 wire \mod.Arithmetic.I_out[72] ;
 wire \mod.Arithmetic.I_out[73] ;
 wire \mod.Arithmetic.I_out[74] ;
 wire \mod.Arithmetic.I_out[75] ;
 wire \mod.Arithmetic.I_out[76] ;
 wire \mod.Arithmetic.I_out[77] ;
 wire \mod.Arithmetic.I_out[78] ;
 wire \mod.Arithmetic.I_out[79] ;
 wire \mod.DM_en ;
 wire \mod.DMen_reg ;
 wire \mod.DMen_reg2 ;
 wire \mod.Data_Mem.F_M.MRAM[0][0] ;
 wire \mod.Data_Mem.F_M.MRAM[0][1] ;
 wire \mod.Data_Mem.F_M.MRAM[0][2] ;
 wire \mod.Data_Mem.F_M.MRAM[0][3] ;
 wire \mod.Data_Mem.F_M.MRAM[0][4] ;
 wire \mod.Data_Mem.F_M.MRAM[0][5] ;
 wire \mod.Data_Mem.F_M.MRAM[0][6] ;
 wire \mod.Data_Mem.F_M.MRAM[0][7] ;
 wire \mod.Data_Mem.F_M.MRAM[10][0] ;
 wire \mod.Data_Mem.F_M.MRAM[10][1] ;
 wire \mod.Data_Mem.F_M.MRAM[10][2] ;
 wire \mod.Data_Mem.F_M.MRAM[10][3] ;
 wire \mod.Data_Mem.F_M.MRAM[10][4] ;
 wire \mod.Data_Mem.F_M.MRAM[10][5] ;
 wire \mod.Data_Mem.F_M.MRAM[10][6] ;
 wire \mod.Data_Mem.F_M.MRAM[10][7] ;
 wire \mod.Data_Mem.F_M.MRAM[11][0] ;
 wire \mod.Data_Mem.F_M.MRAM[11][1] ;
 wire \mod.Data_Mem.F_M.MRAM[11][2] ;
 wire \mod.Data_Mem.F_M.MRAM[11][3] ;
 wire \mod.Data_Mem.F_M.MRAM[11][4] ;
 wire \mod.Data_Mem.F_M.MRAM[11][5] ;
 wire \mod.Data_Mem.F_M.MRAM[11][6] ;
 wire \mod.Data_Mem.F_M.MRAM[11][7] ;
 wire \mod.Data_Mem.F_M.MRAM[12][0] ;
 wire \mod.Data_Mem.F_M.MRAM[12][1] ;
 wire \mod.Data_Mem.F_M.MRAM[12][2] ;
 wire \mod.Data_Mem.F_M.MRAM[12][3] ;
 wire \mod.Data_Mem.F_M.MRAM[12][4] ;
 wire \mod.Data_Mem.F_M.MRAM[12][5] ;
 wire \mod.Data_Mem.F_M.MRAM[12][6] ;
 wire \mod.Data_Mem.F_M.MRAM[12][7] ;
 wire \mod.Data_Mem.F_M.MRAM[13][0] ;
 wire \mod.Data_Mem.F_M.MRAM[13][1] ;
 wire \mod.Data_Mem.F_M.MRAM[13][2] ;
 wire \mod.Data_Mem.F_M.MRAM[13][3] ;
 wire \mod.Data_Mem.F_M.MRAM[13][4] ;
 wire \mod.Data_Mem.F_M.MRAM[13][5] ;
 wire \mod.Data_Mem.F_M.MRAM[13][6] ;
 wire \mod.Data_Mem.F_M.MRAM[13][7] ;
 wire \mod.Data_Mem.F_M.MRAM[14][0] ;
 wire \mod.Data_Mem.F_M.MRAM[14][1] ;
 wire \mod.Data_Mem.F_M.MRAM[14][2] ;
 wire \mod.Data_Mem.F_M.MRAM[14][3] ;
 wire \mod.Data_Mem.F_M.MRAM[14][4] ;
 wire \mod.Data_Mem.F_M.MRAM[14][5] ;
 wire \mod.Data_Mem.F_M.MRAM[14][6] ;
 wire \mod.Data_Mem.F_M.MRAM[14][7] ;
 wire \mod.Data_Mem.F_M.MRAM[15][0] ;
 wire \mod.Data_Mem.F_M.MRAM[15][1] ;
 wire \mod.Data_Mem.F_M.MRAM[15][2] ;
 wire \mod.Data_Mem.F_M.MRAM[15][3] ;
 wire \mod.Data_Mem.F_M.MRAM[15][4] ;
 wire \mod.Data_Mem.F_M.MRAM[15][5] ;
 wire \mod.Data_Mem.F_M.MRAM[15][6] ;
 wire \mod.Data_Mem.F_M.MRAM[15][7] ;
 wire \mod.Data_Mem.F_M.MRAM[16][0] ;
 wire \mod.Data_Mem.F_M.MRAM[16][1] ;
 wire \mod.Data_Mem.F_M.MRAM[16][2] ;
 wire \mod.Data_Mem.F_M.MRAM[16][3] ;
 wire \mod.Data_Mem.F_M.MRAM[16][4] ;
 wire \mod.Data_Mem.F_M.MRAM[16][5] ;
 wire \mod.Data_Mem.F_M.MRAM[16][6] ;
 wire \mod.Data_Mem.F_M.MRAM[16][7] ;
 wire \mod.Data_Mem.F_M.MRAM[17][0] ;
 wire \mod.Data_Mem.F_M.MRAM[17][1] ;
 wire \mod.Data_Mem.F_M.MRAM[17][2] ;
 wire \mod.Data_Mem.F_M.MRAM[17][3] ;
 wire \mod.Data_Mem.F_M.MRAM[17][4] ;
 wire \mod.Data_Mem.F_M.MRAM[17][5] ;
 wire \mod.Data_Mem.F_M.MRAM[17][6] ;
 wire \mod.Data_Mem.F_M.MRAM[17][7] ;
 wire \mod.Data_Mem.F_M.MRAM[18][0] ;
 wire \mod.Data_Mem.F_M.MRAM[18][1] ;
 wire \mod.Data_Mem.F_M.MRAM[18][2] ;
 wire \mod.Data_Mem.F_M.MRAM[18][3] ;
 wire \mod.Data_Mem.F_M.MRAM[18][4] ;
 wire \mod.Data_Mem.F_M.MRAM[18][5] ;
 wire \mod.Data_Mem.F_M.MRAM[18][6] ;
 wire \mod.Data_Mem.F_M.MRAM[18][7] ;
 wire \mod.Data_Mem.F_M.MRAM[19][0] ;
 wire \mod.Data_Mem.F_M.MRAM[19][1] ;
 wire \mod.Data_Mem.F_M.MRAM[19][2] ;
 wire \mod.Data_Mem.F_M.MRAM[19][3] ;
 wire \mod.Data_Mem.F_M.MRAM[19][4] ;
 wire \mod.Data_Mem.F_M.MRAM[19][5] ;
 wire \mod.Data_Mem.F_M.MRAM[19][6] ;
 wire \mod.Data_Mem.F_M.MRAM[19][7] ;
 wire \mod.Data_Mem.F_M.MRAM[1][0] ;
 wire \mod.Data_Mem.F_M.MRAM[1][1] ;
 wire \mod.Data_Mem.F_M.MRAM[1][2] ;
 wire \mod.Data_Mem.F_M.MRAM[1][3] ;
 wire \mod.Data_Mem.F_M.MRAM[1][4] ;
 wire \mod.Data_Mem.F_M.MRAM[1][5] ;
 wire \mod.Data_Mem.F_M.MRAM[1][6] ;
 wire \mod.Data_Mem.F_M.MRAM[1][7] ;
 wire \mod.Data_Mem.F_M.MRAM[20][0] ;
 wire \mod.Data_Mem.F_M.MRAM[20][1] ;
 wire \mod.Data_Mem.F_M.MRAM[20][2] ;
 wire \mod.Data_Mem.F_M.MRAM[20][3] ;
 wire \mod.Data_Mem.F_M.MRAM[20][4] ;
 wire \mod.Data_Mem.F_M.MRAM[20][5] ;
 wire \mod.Data_Mem.F_M.MRAM[20][6] ;
 wire \mod.Data_Mem.F_M.MRAM[20][7] ;
 wire \mod.Data_Mem.F_M.MRAM[21][0] ;
 wire \mod.Data_Mem.F_M.MRAM[21][1] ;
 wire \mod.Data_Mem.F_M.MRAM[21][2] ;
 wire \mod.Data_Mem.F_M.MRAM[21][3] ;
 wire \mod.Data_Mem.F_M.MRAM[21][4] ;
 wire \mod.Data_Mem.F_M.MRAM[21][5] ;
 wire \mod.Data_Mem.F_M.MRAM[21][6] ;
 wire \mod.Data_Mem.F_M.MRAM[21][7] ;
 wire \mod.Data_Mem.F_M.MRAM[22][0] ;
 wire \mod.Data_Mem.F_M.MRAM[22][1] ;
 wire \mod.Data_Mem.F_M.MRAM[22][2] ;
 wire \mod.Data_Mem.F_M.MRAM[22][3] ;
 wire \mod.Data_Mem.F_M.MRAM[22][4] ;
 wire \mod.Data_Mem.F_M.MRAM[22][5] ;
 wire \mod.Data_Mem.F_M.MRAM[22][6] ;
 wire \mod.Data_Mem.F_M.MRAM[22][7] ;
 wire \mod.Data_Mem.F_M.MRAM[23][0] ;
 wire \mod.Data_Mem.F_M.MRAM[23][1] ;
 wire \mod.Data_Mem.F_M.MRAM[23][2] ;
 wire \mod.Data_Mem.F_M.MRAM[23][3] ;
 wire \mod.Data_Mem.F_M.MRAM[23][4] ;
 wire \mod.Data_Mem.F_M.MRAM[23][5] ;
 wire \mod.Data_Mem.F_M.MRAM[23][6] ;
 wire \mod.Data_Mem.F_M.MRAM[23][7] ;
 wire \mod.Data_Mem.F_M.MRAM[24][0] ;
 wire \mod.Data_Mem.F_M.MRAM[24][1] ;
 wire \mod.Data_Mem.F_M.MRAM[24][2] ;
 wire \mod.Data_Mem.F_M.MRAM[24][3] ;
 wire \mod.Data_Mem.F_M.MRAM[24][4] ;
 wire \mod.Data_Mem.F_M.MRAM[24][5] ;
 wire \mod.Data_Mem.F_M.MRAM[24][6] ;
 wire \mod.Data_Mem.F_M.MRAM[24][7] ;
 wire \mod.Data_Mem.F_M.MRAM[25][0] ;
 wire \mod.Data_Mem.F_M.MRAM[25][1] ;
 wire \mod.Data_Mem.F_M.MRAM[25][2] ;
 wire \mod.Data_Mem.F_M.MRAM[25][3] ;
 wire \mod.Data_Mem.F_M.MRAM[25][4] ;
 wire \mod.Data_Mem.F_M.MRAM[25][5] ;
 wire \mod.Data_Mem.F_M.MRAM[25][6] ;
 wire \mod.Data_Mem.F_M.MRAM[25][7] ;
 wire \mod.Data_Mem.F_M.MRAM[26][0] ;
 wire \mod.Data_Mem.F_M.MRAM[26][1] ;
 wire \mod.Data_Mem.F_M.MRAM[26][2] ;
 wire \mod.Data_Mem.F_M.MRAM[26][3] ;
 wire \mod.Data_Mem.F_M.MRAM[26][4] ;
 wire \mod.Data_Mem.F_M.MRAM[26][5] ;
 wire \mod.Data_Mem.F_M.MRAM[26][6] ;
 wire \mod.Data_Mem.F_M.MRAM[26][7] ;
 wire \mod.Data_Mem.F_M.MRAM[27][0] ;
 wire \mod.Data_Mem.F_M.MRAM[27][1] ;
 wire \mod.Data_Mem.F_M.MRAM[27][2] ;
 wire \mod.Data_Mem.F_M.MRAM[27][3] ;
 wire \mod.Data_Mem.F_M.MRAM[27][4] ;
 wire \mod.Data_Mem.F_M.MRAM[27][5] ;
 wire \mod.Data_Mem.F_M.MRAM[27][6] ;
 wire \mod.Data_Mem.F_M.MRAM[27][7] ;
 wire \mod.Data_Mem.F_M.MRAM[28][0] ;
 wire \mod.Data_Mem.F_M.MRAM[28][1] ;
 wire \mod.Data_Mem.F_M.MRAM[28][2] ;
 wire \mod.Data_Mem.F_M.MRAM[28][3] ;
 wire \mod.Data_Mem.F_M.MRAM[28][4] ;
 wire \mod.Data_Mem.F_M.MRAM[28][5] ;
 wire \mod.Data_Mem.F_M.MRAM[28][6] ;
 wire \mod.Data_Mem.F_M.MRAM[28][7] ;
 wire \mod.Data_Mem.F_M.MRAM[29][0] ;
 wire \mod.Data_Mem.F_M.MRAM[29][1] ;
 wire \mod.Data_Mem.F_M.MRAM[29][2] ;
 wire \mod.Data_Mem.F_M.MRAM[29][3] ;
 wire \mod.Data_Mem.F_M.MRAM[29][4] ;
 wire \mod.Data_Mem.F_M.MRAM[29][5] ;
 wire \mod.Data_Mem.F_M.MRAM[29][6] ;
 wire \mod.Data_Mem.F_M.MRAM[29][7] ;
 wire \mod.Data_Mem.F_M.MRAM[2][0] ;
 wire \mod.Data_Mem.F_M.MRAM[2][1] ;
 wire \mod.Data_Mem.F_M.MRAM[2][2] ;
 wire \mod.Data_Mem.F_M.MRAM[2][3] ;
 wire \mod.Data_Mem.F_M.MRAM[2][4] ;
 wire \mod.Data_Mem.F_M.MRAM[2][5] ;
 wire \mod.Data_Mem.F_M.MRAM[2][6] ;
 wire \mod.Data_Mem.F_M.MRAM[2][7] ;
 wire \mod.Data_Mem.F_M.MRAM[30][0] ;
 wire \mod.Data_Mem.F_M.MRAM[30][1] ;
 wire \mod.Data_Mem.F_M.MRAM[30][2] ;
 wire \mod.Data_Mem.F_M.MRAM[30][3] ;
 wire \mod.Data_Mem.F_M.MRAM[30][4] ;
 wire \mod.Data_Mem.F_M.MRAM[30][5] ;
 wire \mod.Data_Mem.F_M.MRAM[30][6] ;
 wire \mod.Data_Mem.F_M.MRAM[30][7] ;
 wire \mod.Data_Mem.F_M.MRAM[31][0] ;
 wire \mod.Data_Mem.F_M.MRAM[31][1] ;
 wire \mod.Data_Mem.F_M.MRAM[31][2] ;
 wire \mod.Data_Mem.F_M.MRAM[31][3] ;
 wire \mod.Data_Mem.F_M.MRAM[31][4] ;
 wire \mod.Data_Mem.F_M.MRAM[31][5] ;
 wire \mod.Data_Mem.F_M.MRAM[31][6] ;
 wire \mod.Data_Mem.F_M.MRAM[31][7] ;
 wire \mod.Data_Mem.F_M.MRAM[3][0] ;
 wire \mod.Data_Mem.F_M.MRAM[3][1] ;
 wire \mod.Data_Mem.F_M.MRAM[3][2] ;
 wire \mod.Data_Mem.F_M.MRAM[3][3] ;
 wire \mod.Data_Mem.F_M.MRAM[3][4] ;
 wire \mod.Data_Mem.F_M.MRAM[3][5] ;
 wire \mod.Data_Mem.F_M.MRAM[3][6] ;
 wire \mod.Data_Mem.F_M.MRAM[3][7] ;
 wire \mod.Data_Mem.F_M.MRAM[4][0] ;
 wire \mod.Data_Mem.F_M.MRAM[4][1] ;
 wire \mod.Data_Mem.F_M.MRAM[4][2] ;
 wire \mod.Data_Mem.F_M.MRAM[4][3] ;
 wire \mod.Data_Mem.F_M.MRAM[4][4] ;
 wire \mod.Data_Mem.F_M.MRAM[4][5] ;
 wire \mod.Data_Mem.F_M.MRAM[4][6] ;
 wire \mod.Data_Mem.F_M.MRAM[4][7] ;
 wire \mod.Data_Mem.F_M.MRAM[5][0] ;
 wire \mod.Data_Mem.F_M.MRAM[5][1] ;
 wire \mod.Data_Mem.F_M.MRAM[5][2] ;
 wire \mod.Data_Mem.F_M.MRAM[5][3] ;
 wire \mod.Data_Mem.F_M.MRAM[5][4] ;
 wire \mod.Data_Mem.F_M.MRAM[5][5] ;
 wire \mod.Data_Mem.F_M.MRAM[5][6] ;
 wire \mod.Data_Mem.F_M.MRAM[5][7] ;
 wire \mod.Data_Mem.F_M.MRAM[6][0] ;
 wire \mod.Data_Mem.F_M.MRAM[6][1] ;
 wire \mod.Data_Mem.F_M.MRAM[6][2] ;
 wire \mod.Data_Mem.F_M.MRAM[6][3] ;
 wire \mod.Data_Mem.F_M.MRAM[6][4] ;
 wire \mod.Data_Mem.F_M.MRAM[6][5] ;
 wire \mod.Data_Mem.F_M.MRAM[6][6] ;
 wire \mod.Data_Mem.F_M.MRAM[6][7] ;
 wire \mod.Data_Mem.F_M.MRAM[768][0] ;
 wire \mod.Data_Mem.F_M.MRAM[768][1] ;
 wire \mod.Data_Mem.F_M.MRAM[768][2] ;
 wire \mod.Data_Mem.F_M.MRAM[768][3] ;
 wire \mod.Data_Mem.F_M.MRAM[768][4] ;
 wire \mod.Data_Mem.F_M.MRAM[768][5] ;
 wire \mod.Data_Mem.F_M.MRAM[768][6] ;
 wire \mod.Data_Mem.F_M.MRAM[768][7] ;
 wire \mod.Data_Mem.F_M.MRAM[769][0] ;
 wire \mod.Data_Mem.F_M.MRAM[769][1] ;
 wire \mod.Data_Mem.F_M.MRAM[769][2] ;
 wire \mod.Data_Mem.F_M.MRAM[769][3] ;
 wire \mod.Data_Mem.F_M.MRAM[769][4] ;
 wire \mod.Data_Mem.F_M.MRAM[769][5] ;
 wire \mod.Data_Mem.F_M.MRAM[769][6] ;
 wire \mod.Data_Mem.F_M.MRAM[769][7] ;
 wire \mod.Data_Mem.F_M.MRAM[770][0] ;
 wire \mod.Data_Mem.F_M.MRAM[770][1] ;
 wire \mod.Data_Mem.F_M.MRAM[770][2] ;
 wire \mod.Data_Mem.F_M.MRAM[770][3] ;
 wire \mod.Data_Mem.F_M.MRAM[770][4] ;
 wire \mod.Data_Mem.F_M.MRAM[770][5] ;
 wire \mod.Data_Mem.F_M.MRAM[770][6] ;
 wire \mod.Data_Mem.F_M.MRAM[770][7] ;
 wire \mod.Data_Mem.F_M.MRAM[771][0] ;
 wire \mod.Data_Mem.F_M.MRAM[771][1] ;
 wire \mod.Data_Mem.F_M.MRAM[771][2] ;
 wire \mod.Data_Mem.F_M.MRAM[771][3] ;
 wire \mod.Data_Mem.F_M.MRAM[771][4] ;
 wire \mod.Data_Mem.F_M.MRAM[771][5] ;
 wire \mod.Data_Mem.F_M.MRAM[771][6] ;
 wire \mod.Data_Mem.F_M.MRAM[771][7] ;
 wire \mod.Data_Mem.F_M.MRAM[772][0] ;
 wire \mod.Data_Mem.F_M.MRAM[772][1] ;
 wire \mod.Data_Mem.F_M.MRAM[772][2] ;
 wire \mod.Data_Mem.F_M.MRAM[772][3] ;
 wire \mod.Data_Mem.F_M.MRAM[772][4] ;
 wire \mod.Data_Mem.F_M.MRAM[772][5] ;
 wire \mod.Data_Mem.F_M.MRAM[772][6] ;
 wire \mod.Data_Mem.F_M.MRAM[772][7] ;
 wire \mod.Data_Mem.F_M.MRAM[773][0] ;
 wire \mod.Data_Mem.F_M.MRAM[773][1] ;
 wire \mod.Data_Mem.F_M.MRAM[773][2] ;
 wire \mod.Data_Mem.F_M.MRAM[773][3] ;
 wire \mod.Data_Mem.F_M.MRAM[773][4] ;
 wire \mod.Data_Mem.F_M.MRAM[773][5] ;
 wire \mod.Data_Mem.F_M.MRAM[773][6] ;
 wire \mod.Data_Mem.F_M.MRAM[773][7] ;
 wire \mod.Data_Mem.F_M.MRAM[774][0] ;
 wire \mod.Data_Mem.F_M.MRAM[774][1] ;
 wire \mod.Data_Mem.F_M.MRAM[774][2] ;
 wire \mod.Data_Mem.F_M.MRAM[774][3] ;
 wire \mod.Data_Mem.F_M.MRAM[774][4] ;
 wire \mod.Data_Mem.F_M.MRAM[774][5] ;
 wire \mod.Data_Mem.F_M.MRAM[774][6] ;
 wire \mod.Data_Mem.F_M.MRAM[774][7] ;
 wire \mod.Data_Mem.F_M.MRAM[775][0] ;
 wire \mod.Data_Mem.F_M.MRAM[775][1] ;
 wire \mod.Data_Mem.F_M.MRAM[775][2] ;
 wire \mod.Data_Mem.F_M.MRAM[775][3] ;
 wire \mod.Data_Mem.F_M.MRAM[775][4] ;
 wire \mod.Data_Mem.F_M.MRAM[775][5] ;
 wire \mod.Data_Mem.F_M.MRAM[775][6] ;
 wire \mod.Data_Mem.F_M.MRAM[775][7] ;
 wire \mod.Data_Mem.F_M.MRAM[776][0] ;
 wire \mod.Data_Mem.F_M.MRAM[776][1] ;
 wire \mod.Data_Mem.F_M.MRAM[776][2] ;
 wire \mod.Data_Mem.F_M.MRAM[776][3] ;
 wire \mod.Data_Mem.F_M.MRAM[776][4] ;
 wire \mod.Data_Mem.F_M.MRAM[776][5] ;
 wire \mod.Data_Mem.F_M.MRAM[776][6] ;
 wire \mod.Data_Mem.F_M.MRAM[776][7] ;
 wire \mod.Data_Mem.F_M.MRAM[777][0] ;
 wire \mod.Data_Mem.F_M.MRAM[777][1] ;
 wire \mod.Data_Mem.F_M.MRAM[777][2] ;
 wire \mod.Data_Mem.F_M.MRAM[777][3] ;
 wire \mod.Data_Mem.F_M.MRAM[777][4] ;
 wire \mod.Data_Mem.F_M.MRAM[777][5] ;
 wire \mod.Data_Mem.F_M.MRAM[777][6] ;
 wire \mod.Data_Mem.F_M.MRAM[777][7] ;
 wire \mod.Data_Mem.F_M.MRAM[778][0] ;
 wire \mod.Data_Mem.F_M.MRAM[778][1] ;
 wire \mod.Data_Mem.F_M.MRAM[778][2] ;
 wire \mod.Data_Mem.F_M.MRAM[778][3] ;
 wire \mod.Data_Mem.F_M.MRAM[778][4] ;
 wire \mod.Data_Mem.F_M.MRAM[778][5] ;
 wire \mod.Data_Mem.F_M.MRAM[778][6] ;
 wire \mod.Data_Mem.F_M.MRAM[778][7] ;
 wire \mod.Data_Mem.F_M.MRAM[779][0] ;
 wire \mod.Data_Mem.F_M.MRAM[779][1] ;
 wire \mod.Data_Mem.F_M.MRAM[779][2] ;
 wire \mod.Data_Mem.F_M.MRAM[779][3] ;
 wire \mod.Data_Mem.F_M.MRAM[779][4] ;
 wire \mod.Data_Mem.F_M.MRAM[779][5] ;
 wire \mod.Data_Mem.F_M.MRAM[779][6] ;
 wire \mod.Data_Mem.F_M.MRAM[779][7] ;
 wire \mod.Data_Mem.F_M.MRAM[780][0] ;
 wire \mod.Data_Mem.F_M.MRAM[780][1] ;
 wire \mod.Data_Mem.F_M.MRAM[780][2] ;
 wire \mod.Data_Mem.F_M.MRAM[780][3] ;
 wire \mod.Data_Mem.F_M.MRAM[780][4] ;
 wire \mod.Data_Mem.F_M.MRAM[780][5] ;
 wire \mod.Data_Mem.F_M.MRAM[780][6] ;
 wire \mod.Data_Mem.F_M.MRAM[780][7] ;
 wire \mod.Data_Mem.F_M.MRAM[781][0] ;
 wire \mod.Data_Mem.F_M.MRAM[781][1] ;
 wire \mod.Data_Mem.F_M.MRAM[781][2] ;
 wire \mod.Data_Mem.F_M.MRAM[781][3] ;
 wire \mod.Data_Mem.F_M.MRAM[781][4] ;
 wire \mod.Data_Mem.F_M.MRAM[781][5] ;
 wire \mod.Data_Mem.F_M.MRAM[781][6] ;
 wire \mod.Data_Mem.F_M.MRAM[781][7] ;
 wire \mod.Data_Mem.F_M.MRAM[782][0] ;
 wire \mod.Data_Mem.F_M.MRAM[782][1] ;
 wire \mod.Data_Mem.F_M.MRAM[782][2] ;
 wire \mod.Data_Mem.F_M.MRAM[782][3] ;
 wire \mod.Data_Mem.F_M.MRAM[782][4] ;
 wire \mod.Data_Mem.F_M.MRAM[782][5] ;
 wire \mod.Data_Mem.F_M.MRAM[782][6] ;
 wire \mod.Data_Mem.F_M.MRAM[782][7] ;
 wire \mod.Data_Mem.F_M.MRAM[783][0] ;
 wire \mod.Data_Mem.F_M.MRAM[783][1] ;
 wire \mod.Data_Mem.F_M.MRAM[783][2] ;
 wire \mod.Data_Mem.F_M.MRAM[783][3] ;
 wire \mod.Data_Mem.F_M.MRAM[783][4] ;
 wire \mod.Data_Mem.F_M.MRAM[783][5] ;
 wire \mod.Data_Mem.F_M.MRAM[783][6] ;
 wire \mod.Data_Mem.F_M.MRAM[783][7] ;
 wire \mod.Data_Mem.F_M.MRAM[784][0] ;
 wire \mod.Data_Mem.F_M.MRAM[784][1] ;
 wire \mod.Data_Mem.F_M.MRAM[784][2] ;
 wire \mod.Data_Mem.F_M.MRAM[784][3] ;
 wire \mod.Data_Mem.F_M.MRAM[784][4] ;
 wire \mod.Data_Mem.F_M.MRAM[784][5] ;
 wire \mod.Data_Mem.F_M.MRAM[784][6] ;
 wire \mod.Data_Mem.F_M.MRAM[784][7] ;
 wire \mod.Data_Mem.F_M.MRAM[785][0] ;
 wire \mod.Data_Mem.F_M.MRAM[785][1] ;
 wire \mod.Data_Mem.F_M.MRAM[785][2] ;
 wire \mod.Data_Mem.F_M.MRAM[785][3] ;
 wire \mod.Data_Mem.F_M.MRAM[785][4] ;
 wire \mod.Data_Mem.F_M.MRAM[785][5] ;
 wire \mod.Data_Mem.F_M.MRAM[785][6] ;
 wire \mod.Data_Mem.F_M.MRAM[785][7] ;
 wire \mod.Data_Mem.F_M.MRAM[786][0] ;
 wire \mod.Data_Mem.F_M.MRAM[786][1] ;
 wire \mod.Data_Mem.F_M.MRAM[786][2] ;
 wire \mod.Data_Mem.F_M.MRAM[786][3] ;
 wire \mod.Data_Mem.F_M.MRAM[786][4] ;
 wire \mod.Data_Mem.F_M.MRAM[786][5] ;
 wire \mod.Data_Mem.F_M.MRAM[786][6] ;
 wire \mod.Data_Mem.F_M.MRAM[786][7] ;
 wire \mod.Data_Mem.F_M.MRAM[787][0] ;
 wire \mod.Data_Mem.F_M.MRAM[787][1] ;
 wire \mod.Data_Mem.F_M.MRAM[787][2] ;
 wire \mod.Data_Mem.F_M.MRAM[787][3] ;
 wire \mod.Data_Mem.F_M.MRAM[787][4] ;
 wire \mod.Data_Mem.F_M.MRAM[787][5] ;
 wire \mod.Data_Mem.F_M.MRAM[787][6] ;
 wire \mod.Data_Mem.F_M.MRAM[787][7] ;
 wire \mod.Data_Mem.F_M.MRAM[788][0] ;
 wire \mod.Data_Mem.F_M.MRAM[788][1] ;
 wire \mod.Data_Mem.F_M.MRAM[788][2] ;
 wire \mod.Data_Mem.F_M.MRAM[788][3] ;
 wire \mod.Data_Mem.F_M.MRAM[788][4] ;
 wire \mod.Data_Mem.F_M.MRAM[788][5] ;
 wire \mod.Data_Mem.F_M.MRAM[788][6] ;
 wire \mod.Data_Mem.F_M.MRAM[788][7] ;
 wire \mod.Data_Mem.F_M.MRAM[789][0] ;
 wire \mod.Data_Mem.F_M.MRAM[789][1] ;
 wire \mod.Data_Mem.F_M.MRAM[789][2] ;
 wire \mod.Data_Mem.F_M.MRAM[789][3] ;
 wire \mod.Data_Mem.F_M.MRAM[789][4] ;
 wire \mod.Data_Mem.F_M.MRAM[789][5] ;
 wire \mod.Data_Mem.F_M.MRAM[789][6] ;
 wire \mod.Data_Mem.F_M.MRAM[789][7] ;
 wire \mod.Data_Mem.F_M.MRAM[790][0] ;
 wire \mod.Data_Mem.F_M.MRAM[790][1] ;
 wire \mod.Data_Mem.F_M.MRAM[790][2] ;
 wire \mod.Data_Mem.F_M.MRAM[790][3] ;
 wire \mod.Data_Mem.F_M.MRAM[790][4] ;
 wire \mod.Data_Mem.F_M.MRAM[790][5] ;
 wire \mod.Data_Mem.F_M.MRAM[790][6] ;
 wire \mod.Data_Mem.F_M.MRAM[790][7] ;
 wire \mod.Data_Mem.F_M.MRAM[791][0] ;
 wire \mod.Data_Mem.F_M.MRAM[791][1] ;
 wire \mod.Data_Mem.F_M.MRAM[791][2] ;
 wire \mod.Data_Mem.F_M.MRAM[791][3] ;
 wire \mod.Data_Mem.F_M.MRAM[791][4] ;
 wire \mod.Data_Mem.F_M.MRAM[791][5] ;
 wire \mod.Data_Mem.F_M.MRAM[791][6] ;
 wire \mod.Data_Mem.F_M.MRAM[791][7] ;
 wire \mod.Data_Mem.F_M.MRAM[792][0] ;
 wire \mod.Data_Mem.F_M.MRAM[792][1] ;
 wire \mod.Data_Mem.F_M.MRAM[792][2] ;
 wire \mod.Data_Mem.F_M.MRAM[792][3] ;
 wire \mod.Data_Mem.F_M.MRAM[792][4] ;
 wire \mod.Data_Mem.F_M.MRAM[792][5] ;
 wire \mod.Data_Mem.F_M.MRAM[792][6] ;
 wire \mod.Data_Mem.F_M.MRAM[792][7] ;
 wire \mod.Data_Mem.F_M.MRAM[793][0] ;
 wire \mod.Data_Mem.F_M.MRAM[793][1] ;
 wire \mod.Data_Mem.F_M.MRAM[793][2] ;
 wire \mod.Data_Mem.F_M.MRAM[793][3] ;
 wire \mod.Data_Mem.F_M.MRAM[793][4] ;
 wire \mod.Data_Mem.F_M.MRAM[793][5] ;
 wire \mod.Data_Mem.F_M.MRAM[793][6] ;
 wire \mod.Data_Mem.F_M.MRAM[793][7] ;
 wire \mod.Data_Mem.F_M.MRAM[794][0] ;
 wire \mod.Data_Mem.F_M.MRAM[794][1] ;
 wire \mod.Data_Mem.F_M.MRAM[794][2] ;
 wire \mod.Data_Mem.F_M.MRAM[794][3] ;
 wire \mod.Data_Mem.F_M.MRAM[794][4] ;
 wire \mod.Data_Mem.F_M.MRAM[794][5] ;
 wire \mod.Data_Mem.F_M.MRAM[794][6] ;
 wire \mod.Data_Mem.F_M.MRAM[794][7] ;
 wire \mod.Data_Mem.F_M.MRAM[795][0] ;
 wire \mod.Data_Mem.F_M.MRAM[795][1] ;
 wire \mod.Data_Mem.F_M.MRAM[795][2] ;
 wire \mod.Data_Mem.F_M.MRAM[795][3] ;
 wire \mod.Data_Mem.F_M.MRAM[795][4] ;
 wire \mod.Data_Mem.F_M.MRAM[795][5] ;
 wire \mod.Data_Mem.F_M.MRAM[795][6] ;
 wire \mod.Data_Mem.F_M.MRAM[795][7] ;
 wire \mod.Data_Mem.F_M.MRAM[796][0] ;
 wire \mod.Data_Mem.F_M.MRAM[796][1] ;
 wire \mod.Data_Mem.F_M.MRAM[796][2] ;
 wire \mod.Data_Mem.F_M.MRAM[796][3] ;
 wire \mod.Data_Mem.F_M.MRAM[796][4] ;
 wire \mod.Data_Mem.F_M.MRAM[796][5] ;
 wire \mod.Data_Mem.F_M.MRAM[796][6] ;
 wire \mod.Data_Mem.F_M.MRAM[796][7] ;
 wire \mod.Data_Mem.F_M.MRAM[797][0] ;
 wire \mod.Data_Mem.F_M.MRAM[797][1] ;
 wire \mod.Data_Mem.F_M.MRAM[797][2] ;
 wire \mod.Data_Mem.F_M.MRAM[797][3] ;
 wire \mod.Data_Mem.F_M.MRAM[797][4] ;
 wire \mod.Data_Mem.F_M.MRAM[797][5] ;
 wire \mod.Data_Mem.F_M.MRAM[797][6] ;
 wire \mod.Data_Mem.F_M.MRAM[797][7] ;
 wire \mod.Data_Mem.F_M.MRAM[798][0] ;
 wire \mod.Data_Mem.F_M.MRAM[798][1] ;
 wire \mod.Data_Mem.F_M.MRAM[798][2] ;
 wire \mod.Data_Mem.F_M.MRAM[798][3] ;
 wire \mod.Data_Mem.F_M.MRAM[798][4] ;
 wire \mod.Data_Mem.F_M.MRAM[798][5] ;
 wire \mod.Data_Mem.F_M.MRAM[798][6] ;
 wire \mod.Data_Mem.F_M.MRAM[798][7] ;
 wire \mod.Data_Mem.F_M.MRAM[799][0] ;
 wire \mod.Data_Mem.F_M.MRAM[799][1] ;
 wire \mod.Data_Mem.F_M.MRAM[799][2] ;
 wire \mod.Data_Mem.F_M.MRAM[799][3] ;
 wire \mod.Data_Mem.F_M.MRAM[799][4] ;
 wire \mod.Data_Mem.F_M.MRAM[799][5] ;
 wire \mod.Data_Mem.F_M.MRAM[799][6] ;
 wire \mod.Data_Mem.F_M.MRAM[799][7] ;
 wire \mod.Data_Mem.F_M.MRAM[7][0] ;
 wire \mod.Data_Mem.F_M.MRAM[7][1] ;
 wire \mod.Data_Mem.F_M.MRAM[7][2] ;
 wire \mod.Data_Mem.F_M.MRAM[7][3] ;
 wire \mod.Data_Mem.F_M.MRAM[7][4] ;
 wire \mod.Data_Mem.F_M.MRAM[7][5] ;
 wire \mod.Data_Mem.F_M.MRAM[7][6] ;
 wire \mod.Data_Mem.F_M.MRAM[7][7] ;
 wire \mod.Data_Mem.F_M.MRAM[8][0] ;
 wire \mod.Data_Mem.F_M.MRAM[8][1] ;
 wire \mod.Data_Mem.F_M.MRAM[8][2] ;
 wire \mod.Data_Mem.F_M.MRAM[8][3] ;
 wire \mod.Data_Mem.F_M.MRAM[8][4] ;
 wire \mod.Data_Mem.F_M.MRAM[8][5] ;
 wire \mod.Data_Mem.F_M.MRAM[8][6] ;
 wire \mod.Data_Mem.F_M.MRAM[8][7] ;
 wire \mod.Data_Mem.F_M.MRAM[9][0] ;
 wire \mod.Data_Mem.F_M.MRAM[9][1] ;
 wire \mod.Data_Mem.F_M.MRAM[9][2] ;
 wire \mod.Data_Mem.F_M.MRAM[9][3] ;
 wire \mod.Data_Mem.F_M.MRAM[9][4] ;
 wire \mod.Data_Mem.F_M.MRAM[9][5] ;
 wire \mod.Data_Mem.F_M.MRAM[9][6] ;
 wire \mod.Data_Mem.F_M.MRAM[9][7] ;
 wire \mod.Data_Mem.F_M.dest[0] ;
 wire \mod.Data_Mem.F_M.dest[1] ;
 wire \mod.Data_Mem.F_M.dest[2] ;
 wire \mod.Data_Mem.F_M.dest[4] ;
 wire \mod.Data_Mem.F_M.dest[8] ;
 wire \mod.Data_Mem.F_M.out_data[0] ;
 wire \mod.Data_Mem.F_M.out_data[10] ;
 wire \mod.Data_Mem.F_M.out_data[11] ;
 wire \mod.Data_Mem.F_M.out_data[12] ;
 wire \mod.Data_Mem.F_M.out_data[13] ;
 wire \mod.Data_Mem.F_M.out_data[14] ;
 wire \mod.Data_Mem.F_M.out_data[15] ;
 wire \mod.Data_Mem.F_M.out_data[16] ;
 wire \mod.Data_Mem.F_M.out_data[17] ;
 wire \mod.Data_Mem.F_M.out_data[18] ;
 wire \mod.Data_Mem.F_M.out_data[19] ;
 wire \mod.Data_Mem.F_M.out_data[1] ;
 wire \mod.Data_Mem.F_M.out_data[20] ;
 wire \mod.Data_Mem.F_M.out_data[21] ;
 wire \mod.Data_Mem.F_M.out_data[22] ;
 wire \mod.Data_Mem.F_M.out_data[23] ;
 wire \mod.Data_Mem.F_M.out_data[24] ;
 wire \mod.Data_Mem.F_M.out_data[25] ;
 wire \mod.Data_Mem.F_M.out_data[26] ;
 wire \mod.Data_Mem.F_M.out_data[27] ;
 wire \mod.Data_Mem.F_M.out_data[28] ;
 wire \mod.Data_Mem.F_M.out_data[29] ;
 wire \mod.Data_Mem.F_M.out_data[2] ;
 wire \mod.Data_Mem.F_M.out_data[30] ;
 wire \mod.Data_Mem.F_M.out_data[31] ;
 wire \mod.Data_Mem.F_M.out_data[32] ;
 wire \mod.Data_Mem.F_M.out_data[33] ;
 wire \mod.Data_Mem.F_M.out_data[34] ;
 wire \mod.Data_Mem.F_M.out_data[35] ;
 wire \mod.Data_Mem.F_M.out_data[36] ;
 wire \mod.Data_Mem.F_M.out_data[37] ;
 wire \mod.Data_Mem.F_M.out_data[38] ;
 wire \mod.Data_Mem.F_M.out_data[39] ;
 wire \mod.Data_Mem.F_M.out_data[3] ;
 wire \mod.Data_Mem.F_M.out_data[40] ;
 wire \mod.Data_Mem.F_M.out_data[41] ;
 wire \mod.Data_Mem.F_M.out_data[42] ;
 wire \mod.Data_Mem.F_M.out_data[43] ;
 wire \mod.Data_Mem.F_M.out_data[44] ;
 wire \mod.Data_Mem.F_M.out_data[45] ;
 wire \mod.Data_Mem.F_M.out_data[46] ;
 wire \mod.Data_Mem.F_M.out_data[47] ;
 wire \mod.Data_Mem.F_M.out_data[48] ;
 wire \mod.Data_Mem.F_M.out_data[49] ;
 wire \mod.Data_Mem.F_M.out_data[4] ;
 wire \mod.Data_Mem.F_M.out_data[50] ;
 wire \mod.Data_Mem.F_M.out_data[51] ;
 wire \mod.Data_Mem.F_M.out_data[52] ;
 wire \mod.Data_Mem.F_M.out_data[53] ;
 wire \mod.Data_Mem.F_M.out_data[54] ;
 wire \mod.Data_Mem.F_M.out_data[55] ;
 wire \mod.Data_Mem.F_M.out_data[56] ;
 wire \mod.Data_Mem.F_M.out_data[57] ;
 wire \mod.Data_Mem.F_M.out_data[58] ;
 wire \mod.Data_Mem.F_M.out_data[59] ;
 wire \mod.Data_Mem.F_M.out_data[5] ;
 wire \mod.Data_Mem.F_M.out_data[60] ;
 wire \mod.Data_Mem.F_M.out_data[61] ;
 wire \mod.Data_Mem.F_M.out_data[62] ;
 wire \mod.Data_Mem.F_M.out_data[63] ;
 wire \mod.Data_Mem.F_M.out_data[64] ;
 wire \mod.Data_Mem.F_M.out_data[65] ;
 wire \mod.Data_Mem.F_M.out_data[66] ;
 wire \mod.Data_Mem.F_M.out_data[67] ;
 wire \mod.Data_Mem.F_M.out_data[68] ;
 wire \mod.Data_Mem.F_M.out_data[69] ;
 wire \mod.Data_Mem.F_M.out_data[6] ;
 wire \mod.Data_Mem.F_M.out_data[70] ;
 wire \mod.Data_Mem.F_M.out_data[71] ;
 wire \mod.Data_Mem.F_M.out_data[72] ;
 wire \mod.Data_Mem.F_M.out_data[73] ;
 wire \mod.Data_Mem.F_M.out_data[74] ;
 wire \mod.Data_Mem.F_M.out_data[75] ;
 wire \mod.Data_Mem.F_M.out_data[76] ;
 wire \mod.Data_Mem.F_M.out_data[77] ;
 wire \mod.Data_Mem.F_M.out_data[78] ;
 wire \mod.Data_Mem.F_M.out_data[79] ;
 wire \mod.Data_Mem.F_M.out_data[7] ;
 wire \mod.Data_Mem.F_M.out_data[8] ;
 wire \mod.Data_Mem.F_M.out_data[9] ;
 wire \mod.Data_Mem.F_M.src[0] ;
 wire \mod.Data_Mem.F_M.src[1] ;
 wire \mod.Data_Mem.F_M.src[2] ;
 wire \mod.Data_Mem.F_M.src[4] ;
 wire \mod.Data_Mem.F_M.src[8] ;
 wire \mod.I_addr[0] ;
 wire \mod.I_addr[1] ;
 wire \mod.I_addr[2] ;
 wire \mod.I_addr[3] ;
 wire \mod.I_addr[4] ;
 wire \mod.I_addr[5] ;
 wire \mod.I_addr[6] ;
 wire \mod.I_addr[7] ;
 wire \mod.Instr_Mem.instruction[10] ;
 wire \mod.Instr_Mem.instruction[11] ;
 wire \mod.Instr_Mem.instruction[13] ;
 wire \mod.Instr_Mem.instruction[17] ;
 wire \mod.Instr_Mem.instruction[22] ;
 wire \mod.Instr_Mem.instruction[23] ;
 wire \mod.Instr_Mem.instruction[24] ;
 wire \mod.Instr_Mem.instruction[26] ;
 wire \mod.Instr_Mem.instruction[30] ;
 wire \mod.Instr_Mem.instruction[7] ;
 wire \mod.Instr_Mem.instruction[8] ;
 wire \mod.Instr_Mem.instruction[9] ;
 wire \mod.P1.instr_reg[10] ;
 wire \mod.P1.instr_reg[11] ;
 wire \mod.P1.instr_reg[13] ;
 wire \mod.P1.instr_reg[17] ;
 wire \mod.P1.instr_reg[7] ;
 wire \mod.P1.instr_reg[8] ;
 wire \mod.P1.instr_reg[9] ;
 wire \mod.P2.Rout_reg1[0] ;
 wire \mod.P2.Rout_reg1[1] ;
 wire \mod.P2.Rout_reg[0] ;
 wire \mod.P2.Rout_reg[1] ;
 wire \mod.P2.dest_reg1[0] ;
 wire \mod.P2.dest_reg1[1] ;
 wire \mod.P2.dest_reg1[2] ;
 wire \mod.P2.dest_reg1[4] ;
 wire \mod.P2.dest_reg1[8] ;
 wire \mod.P2.dest_reg[0] ;
 wire \mod.P2.dest_reg[1] ;
 wire \mod.P2.dest_reg[2] ;
 wire \mod.P2.dest_reg[4] ;
 wire \mod.P2.dest_reg[8] ;
 wire \mod.P3.Res[0] ;
 wire \mod.P3.Res[1] ;
 wire \mod.P3.Res[2] ;
 wire \mod.P3.Res[3] ;
 wire \mod.P3.Res[4] ;
 wire \mod.P3.Res[5] ;
 wire \mod.P3.Res[6] ;
 wire \mod.P3.Res[7] ;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net532;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net533;
 wire net561;
 wire net562;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;

 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3933_ (.I(\mod.I_addr[0] ),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3934_ (.I(_0612_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3935_ (.I(\mod.Arithmetic.CN.F_in[0] ),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3936_ (.I(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3937_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3938_ (.I(_0615_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3939_ (.I(_0616_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3940_ (.I(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3941_ (.I(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3942_ (.I(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3943_ (.I(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3944_ (.I(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3945_ (.I(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3946_ (.I(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3947_ (.I(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3948_ (.A1(\mod.P1.instr_reg[17] ),
    .A2(_0625_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3949_ (.I(_0626_),
    .Z(\mod.DM_en ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3950_ (.A1(\mod.P2.Rout_reg[0] ),
    .A2(\mod.P2.Rout_reg[1] ),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3951_ (.I(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3952_ (.I(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3953_ (.I(\mod.Arithmetic.CN.I_in[8] ),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3954_ (.A1(_0623_),
    .A2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3955_ (.I(_0614_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3956_ (.I(_0632_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3957_ (.I(_0633_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3958_ (.I(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3959_ (.I(_0635_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3960_ (.I(\mod.Arithmetic.CN.I_in[16] ),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3961_ (.A1(_0636_),
    .A2(\mod.Arithmetic.CN.I_in[24] ),
    .A3(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3962_ (.I(\mod.Arithmetic.CN.F_in[0] ),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3963_ (.I(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3964_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3965_ (.I(_0641_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3966_ (.I(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3967_ (.I(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3968_ (.A1(_0644_),
    .A2(\mod.Arithmetic.CN.I_in[16] ),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3969_ (.I(_0639_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3970_ (.I(_0646_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3971_ (.I(_0647_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3972_ (.I(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3973_ (.A1(_0649_),
    .A2(\mod.Arithmetic.CN.I_in[24] ),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3974_ (.A1(_0645_),
    .A2(_0650_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3975_ (.A1(_0638_),
    .A2(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3976_ (.A1(_0631_),
    .A2(_0652_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3977_ (.A1(_0619_),
    .A2(\mod.Arithmetic.CN.I_in[32] ),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3978_ (.I(_0635_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3979_ (.I(\mod.Arithmetic.CN.I_in[40] ),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3980_ (.A1(_0655_),
    .A2(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3981_ (.I(_0649_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3982_ (.I(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3983_ (.A1(_0659_),
    .A2(\mod.Arithmetic.CN.I_in[48] ),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3984_ (.I(_0616_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3985_ (.A1(_0661_),
    .A2(\mod.Arithmetic.CN.I_in[56] ),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3986_ (.I(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3987_ (.I(_0661_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3988_ (.I(\mod.Arithmetic.ACTI.x[0] ),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3989_ (.A1(_0664_),
    .A2(_0665_),
    .A3(\mod.Arithmetic.CN.I_in[64] ),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3990_ (.I(\mod.Arithmetic.CN.F_in[0] ),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3991_ (.I(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3992_ (.A1(_0668_),
    .A2(\mod.Arithmetic.CN.I_in[64] ),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3993_ (.A1(_0632_),
    .A2(\mod.Arithmetic.ACTI.x[0] ),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3994_ (.I(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3995_ (.A1(_0669_),
    .A2(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3996_ (.A1(_0666_),
    .A2(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3997_ (.A1(_0663_),
    .A2(_0673_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3998_ (.A1(_0660_),
    .A2(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3999_ (.A1(_0654_),
    .A2(_0657_),
    .A3(_0675_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4000_ (.A1(_0653_),
    .A2(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4001_ (.I(\mod.P2.Rout_reg[1] ),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4002_ (.I(\mod.Arithmetic.ACTI.x[7] ),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4003_ (.I(\mod.Arithmetic.CN.I_in[23] ),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4004_ (.I(\mod.Arithmetic.CN.I_in[15] ),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4005_ (.A1(_0680_),
    .A2(\mod.Arithmetic.I_out[79] ),
    .A3(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4006_ (.I(\mod.Arithmetic.I_out[79] ),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4007_ (.I(\mod.Arithmetic.CN.I_in[21] ),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4008_ (.I(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4009_ (.I(\mod.Arithmetic.CN.I_in[19] ),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4010_ (.I(\mod.Arithmetic.I_out[75] ),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4011_ (.I(\mod.Arithmetic.CN.I_in[18] ),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4012_ (.I(\mod.Arithmetic.I_out[74] ),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4013_ (.I(\mod.Arithmetic.CN.I_in[17] ),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4014_ (.I(_0637_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4015_ (.A1(_0690_),
    .A2(\mod.Arithmetic.I_out[73] ),
    .B(\mod.Arithmetic.I_out[72] ),
    .C(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4016_ (.I(_0688_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4017_ (.A1(_0693_),
    .A2(\mod.Arithmetic.I_out[74] ),
    .B1(_0690_),
    .B2(\mod.Arithmetic.I_out[73] ),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_4 _4018_ (.A1(_0686_),
    .A2(_0687_),
    .B1(_0688_),
    .B2(_0689_),
    .C1(_0692_),
    .C2(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4019_ (.I(\mod.Arithmetic.I_out[76] ),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4020_ (.I(\mod.Arithmetic.CN.I_in[20] ),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4021_ (.A1(_0696_),
    .A2(_0697_),
    .B1(_0686_),
    .B2(_0687_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4022_ (.A1(_0696_),
    .A2(_0697_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4023_ (.A1(_0685_),
    .A2(\mod.Arithmetic.I_out[77] ),
    .B1(_0695_),
    .B2(_0698_),
    .C(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4024_ (.I(\mod.Arithmetic.CN.I_in[22] ),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4025_ (.I(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4026_ (.A1(\mod.Arithmetic.CN.I_in[23] ),
    .A2(_0683_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4027_ (.I(\mod.Arithmetic.I_out[77] ),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4028_ (.A1(_0702_),
    .A2(\mod.Arithmetic.I_out[78] ),
    .B1(_0684_),
    .B2(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4029_ (.A1(_0702_),
    .A2(\mod.Arithmetic.I_out[78] ),
    .B(_0703_),
    .C(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4030_ (.A1(_0702_),
    .A2(\mod.Arithmetic.I_out[78] ),
    .A3(_0703_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4031_ (.A1(\mod.Arithmetic.CN.I_in[23] ),
    .A2(_0683_),
    .B1(_0700_),
    .B2(_0706_),
    .C(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4032_ (.I(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4033_ (.I0(_0637_),
    .I1(\mod.Arithmetic.I_out[72] ),
    .S(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4034_ (.A1(_0680_),
    .A2(\mod.Arithmetic.I_out[79] ),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4035_ (.A1(_0681_),
    .A2(_0711_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4036_ (.I(\mod.Arithmetic.CN.I_in[10] ),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4037_ (.I0(_0688_),
    .I1(\mod.Arithmetic.I_out[74] ),
    .S(_0709_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4038_ (.I(\mod.Arithmetic.CN.I_in[9] ),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4039_ (.I(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4040_ (.I(\mod.Arithmetic.I_out[73] ),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4041_ (.I0(_0690_),
    .I1(_0717_),
    .S(_0708_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4042_ (.I(_0708_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4043_ (.I0(_0693_),
    .I1(_0689_),
    .S(_0719_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4044_ (.I(\mod.Arithmetic.CN.I_in[10] ),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4045_ (.I(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4046_ (.A1(_0716_),
    .A2(_0718_),
    .B1(_0720_),
    .B2(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4047_ (.I(\mod.Arithmetic.I_out[72] ),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4048_ (.I0(_0691_),
    .I1(_0724_),
    .S(_0708_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4049_ (.A1(_0716_),
    .A2(_0718_),
    .B(_0725_),
    .C(_0630_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4050_ (.I0(_0686_),
    .I1(\mod.Arithmetic.I_out[75] ),
    .S(_0719_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4051_ (.I(\mod.Arithmetic.CN.I_in[11] ),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _4052_ (.A1(_0713_),
    .A2(_0714_),
    .B1(_0723_),
    .B2(_0726_),
    .C1(_0727_),
    .C2(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4053_ (.I(\mod.Arithmetic.CN.I_in[12] ),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4054_ (.I(_0730_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4055_ (.I(_0697_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4056_ (.I0(_0732_),
    .I1(_0696_),
    .S(_0719_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4057_ (.A1(_0731_),
    .A2(_0733_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4058_ (.A1(_0728_),
    .A2(_0727_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4059_ (.I0(_0685_),
    .I1(_0704_),
    .S(_0719_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4060_ (.I(\mod.Arithmetic.CN.I_in[13] ),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4061_ (.I(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4062_ (.A1(_0731_),
    .A2(_0733_),
    .B1(_0736_),
    .B2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4063_ (.I(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4064_ (.A1(_0729_),
    .A2(_0734_),
    .A3(_0735_),
    .B(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4065_ (.A1(_0738_),
    .A2(_0736_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4066_ (.I(\mod.Arithmetic.CN.I_in[14] ),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4067_ (.I(_0743_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4068_ (.A1(_0680_),
    .A2(_0683_),
    .B1(_0700_),
    .B2(_0706_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4069_ (.I(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4070_ (.A1(\mod.Arithmetic.I_out[78] ),
    .A2(_0746_),
    .B1(_0709_),
    .B2(\mod.Arithmetic.CN.I_in[22] ),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4071_ (.A1(_0744_),
    .A2(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4072_ (.A1(_0742_),
    .A2(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4073_ (.A1(\mod.Arithmetic.CN.I_in[15] ),
    .A2(_0711_),
    .B1(_0747_),
    .B2(_0744_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4074_ (.A1(_0741_),
    .A2(_0749_),
    .B(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4075_ (.A1(_0712_),
    .A2(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4076_ (.I0(_0630_),
    .I1(_0710_),
    .S(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4077_ (.I(\mod.Arithmetic.ACTI.x[1] ),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4078_ (.A1(_0681_),
    .A2(_0711_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4079_ (.I(_0716_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4080_ (.I0(\mod.Arithmetic.CN.I_in[17] ),
    .I1(\mod.Arithmetic.I_out[73] ),
    .S(_0709_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4081_ (.I(_0630_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4082_ (.A1(_0756_),
    .A2(_0757_),
    .B(_0710_),
    .C(_0758_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4083_ (.I(_0713_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4084_ (.A1(_0756_),
    .A2(_0757_),
    .B1(_0714_),
    .B2(_0760_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4085_ (.A1(_0760_),
    .A2(_0714_),
    .B1(_0727_),
    .B2(_0728_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4086_ (.A1(_0759_),
    .A2(_0761_),
    .B(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4087_ (.A1(_0734_),
    .A2(_0735_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4088_ (.A1(_0763_),
    .A2(_0764_),
    .B(_0739_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4089_ (.A1(_0742_),
    .A2(_0748_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4090_ (.I(_0750_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4091_ (.A1(_0765_),
    .A2(_0766_),
    .B(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4092_ (.A1(_0755_),
    .A2(_0768_),
    .B(_0716_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4093_ (.A1(_0712_),
    .A2(_0757_),
    .A3(_0751_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4094_ (.A1(_0754_),
    .A2(_0769_),
    .A3(_0770_),
    .B(_0665_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4095_ (.I(_0752_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4096_ (.A1(_0755_),
    .A2(_0714_),
    .A3(_0768_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4097_ (.I(\mod.Arithmetic.ACTI.x[2] ),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4098_ (.A1(_0760_),
    .A2(_0772_),
    .B(_0773_),
    .C(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4099_ (.A1(_0769_),
    .A2(_0770_),
    .B(_0754_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4100_ (.A1(_0753_),
    .A2(_0771_),
    .B(_0775_),
    .C(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4101_ (.I(_0774_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4102_ (.A1(_0760_),
    .A2(_0772_),
    .B(_0773_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4103_ (.I0(\mod.Arithmetic.CN.I_in[11] ),
    .I1(_0727_),
    .S(_0752_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4104_ (.I(\mod.Arithmetic.ACTI.x[3] ),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4105_ (.I(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4106_ (.A1(_0778_),
    .A2(_0779_),
    .B1(_0780_),
    .B2(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4107_ (.I(_0752_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4108_ (.A1(_0733_),
    .A2(_0772_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4109_ (.A1(_0731_),
    .A2(_0784_),
    .B(_0785_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4110_ (.I(\mod.Arithmetic.ACTI.x[4] ),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4111_ (.A1(_0782_),
    .A2(_0780_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4112_ (.A1(_0777_),
    .A2(_0783_),
    .B1(_0786_),
    .B2(_0787_),
    .C(_0788_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4113_ (.A1(_0736_),
    .A2(_0784_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4114_ (.A1(_0738_),
    .A2(_0784_),
    .B(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4115_ (.I(\mod.Arithmetic.ACTI.x[5] ),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4116_ (.A1(_0787_),
    .A2(_0786_),
    .B1(_0791_),
    .B2(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4117_ (.A1(_0747_),
    .A2(_0772_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4118_ (.A1(_0744_),
    .A2(_0784_),
    .B(_0794_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4119_ (.A1(_0792_),
    .A2(_0791_),
    .B1(_0795_),
    .B2(\mod.Arithmetic.ACTI.x[6] ),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4120_ (.A1(_0789_),
    .A2(_0793_),
    .B(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4121_ (.A1(\mod.Arithmetic.ACTI.x[7] ),
    .A2(_0682_),
    .B1(_0795_),
    .B2(\mod.Arithmetic.ACTI.x[6] ),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4122_ (.I(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4123_ (.A1(_0679_),
    .A2(_0682_),
    .B1(_0797_),
    .B2(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4124_ (.I(_0800_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4125_ (.A1(_0678_),
    .A2(_0679_),
    .B1(_0801_),
    .B2(\mod.P2.Rout_reg[0] ),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4126_ (.I(\mod.P2.Rout_reg[0] ),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4127_ (.A1(_0803_),
    .A2(_0753_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4128_ (.I(_0801_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4129_ (.A1(_0665_),
    .A2(_0802_),
    .B1(_0804_),
    .B2(_0805_),
    .C(_0628_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4130_ (.A1(_0629_),
    .A2(_0677_),
    .B(_0806_),
    .ZN(\mod.P3.Res[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4131_ (.A1(_0653_),
    .A2(_0676_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4132_ (.A1(_0631_),
    .A2(_0652_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4133_ (.A1(_0632_),
    .A2(\mod.Arithmetic.CN.I_in[17] ),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4134_ (.I(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4135_ (.I(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4136_ (.A1(_0615_),
    .A2(\mod.Arithmetic.CN.I_in[25] ),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4137_ (.I(_0812_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4138_ (.A1(_0650_),
    .A2(_0813_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4139_ (.A1(_0645_),
    .A2(_0811_),
    .A3(_0814_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4140_ (.A1(_0638_),
    .A2(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4141_ (.I(_0636_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4142_ (.A1(_0817_),
    .A2(_0715_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4143_ (.A1(_0631_),
    .A2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4144_ (.A1(_0621_),
    .A2(\mod.Arithmetic.CN.I_in[8] ),
    .A3(_0715_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4145_ (.A1(_0819_),
    .A2(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4146_ (.A1(_0816_),
    .A2(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4147_ (.A1(_0808_),
    .A2(_0822_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4148_ (.I(\mod.Arithmetic.CN.I_in[32] ),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4149_ (.A1(_0621_),
    .A2(_0656_),
    .A3(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4150_ (.A1(_0654_),
    .A2(_0657_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4151_ (.A1(_0825_),
    .A2(_0826_),
    .A3(_0675_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4152_ (.I(_0817_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4153_ (.A1(_0828_),
    .A2(\mod.Arithmetic.CN.I_in[48] ),
    .A3(_0674_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4154_ (.A1(_0635_),
    .A2(\mod.Arithmetic.CN.I_in[33] ),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4155_ (.A1(_0654_),
    .A2(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4156_ (.A1(_0655_),
    .A2(_0824_),
    .A3(\mod.Arithmetic.CN.I_in[33] ),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4157_ (.A1(_0831_),
    .A2(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4158_ (.I(_0618_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4159_ (.A1(_0834_),
    .A2(\mod.Arithmetic.CN.I_in[41] ),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4160_ (.A1(_0657_),
    .A2(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4161_ (.A1(_0659_),
    .A2(\mod.Arithmetic.CN.I_in[40] ),
    .A3(\mod.Arithmetic.CN.I_in[41] ),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4162_ (.A1(_0836_),
    .A2(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4163_ (.A1(_0833_),
    .A2(_0838_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4164_ (.A1(_0825_),
    .A2(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4165_ (.A1(_0663_),
    .A2(_0673_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4166_ (.A1(_0617_),
    .A2(\mod.Arithmetic.CN.I_in[49] ),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4167_ (.A1(_0660_),
    .A2(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4168_ (.A1(_0617_),
    .A2(\mod.Arithmetic.CN.I_in[57] ),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4169_ (.A1(_0662_),
    .A2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4170_ (.A1(_0668_),
    .A2(\mod.Arithmetic.CN.I_in[65] ),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4171_ (.A1(_0668_),
    .A2(\mod.Arithmetic.ACTI.x[1] ),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4172_ (.A1(_0669_),
    .A2(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4173_ (.A1(_0671_),
    .A2(_0846_),
    .A3(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4174_ (.A1(_0666_),
    .A2(_0845_),
    .A3(_0849_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4175_ (.A1(_0841_),
    .A2(_0843_),
    .A3(_0850_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4176_ (.A1(_0829_),
    .A2(_0840_),
    .A3(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4177_ (.A1(_0827_),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4178_ (.A1(_0823_),
    .A2(_0853_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4179_ (.A1(_0807_),
    .A2(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4180_ (.A1(_0678_),
    .A2(_0679_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4181_ (.I(_0856_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4182_ (.A1(_0803_),
    .A2(\mod.P2.Rout_reg[1] ),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4183_ (.I(_0858_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4184_ (.A1(_0769_),
    .A2(_0770_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4185_ (.I0(_0754_),
    .I1(_0860_),
    .S(_0800_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4186_ (.A1(_0754_),
    .A2(_0857_),
    .B1(_0859_),
    .B2(_0861_),
    .C(_0628_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4187_ (.A1(_0629_),
    .A2(_0855_),
    .B(_0862_),
    .ZN(\mod.P3.Res[1] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4188_ (.A1(_0807_),
    .A2(_0854_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4189_ (.A1(_0808_),
    .A2(_0822_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4190_ (.A1(_0825_),
    .A2(_0826_),
    .A3(_0675_),
    .A4(_0852_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4191_ (.A1(_0823_),
    .A2(_0853_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4192_ (.A1(_0865_),
    .A2(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4193_ (.A1(_0816_),
    .A2(_0821_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4194_ (.A1(_0623_),
    .A2(_0656_),
    .A3(_0824_),
    .A4(_0839_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4195_ (.A1(_0638_),
    .A2(_0815_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4196_ (.A1(_0645_),
    .A2(_0810_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4197_ (.A1(_0637_),
    .A2(_0811_),
    .B1(_0871_),
    .B2(_0814_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4198_ (.I(\mod.Arithmetic.CN.I_in[26] ),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4199_ (.A1(\mod.Arithmetic.CN.I_in[24] ),
    .A2(_0873_),
    .A3(_0812_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4200_ (.A1(_0615_),
    .A2(_0873_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4201_ (.A1(\mod.Arithmetic.CN.I_in[24] ),
    .A2(_0813_),
    .B(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4202_ (.A1(_0641_),
    .A2(\mod.Arithmetic.CN.I_in[18] ),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4203_ (.A1(_0809_),
    .A2(_0877_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4204_ (.A1(_0874_),
    .A2(_0876_),
    .B(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4205_ (.I(_0879_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4206_ (.A1(_0878_),
    .A2(_0874_),
    .A3(_0876_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4207_ (.A1(_0880_),
    .A2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4208_ (.A1(_0870_),
    .A2(_0872_),
    .A3(_0882_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4209_ (.A1(_0817_),
    .A2(_0721_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4210_ (.A1(\mod.Arithmetic.CN.I_in[8] ),
    .A2(_0818_),
    .B(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4211_ (.A1(\mod.Arithmetic.CN.I_in[8] ),
    .A2(_0713_),
    .A3(_0818_),
    .B(_0885_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4212_ (.A1(_0883_),
    .A2(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4213_ (.A1(_0869_),
    .A2(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4214_ (.A1(_0829_),
    .A2(_0851_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4215_ (.A1(_0829_),
    .A2(_0851_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4216_ (.A1(_0840_),
    .A2(_0889_),
    .B(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4217_ (.A1(_0833_),
    .A2(_0838_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4218_ (.A1(_0644_),
    .A2(\mod.Arithmetic.CN.I_in[34] ),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4219_ (.I(\mod.Arithmetic.CN.I_in[34] ),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4220_ (.A1(_0824_),
    .A2(_0830_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4221_ (.I0(_0893_),
    .I1(_0894_),
    .S(_0895_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4222_ (.A1(_0634_),
    .A2(\mod.Arithmetic.CN.I_in[42] ),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4223_ (.I(\mod.Arithmetic.CN.I_in[42] ),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4224_ (.A1(_0656_),
    .A2(_0835_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4225_ (.I0(_0897_),
    .I1(_0898_),
    .S(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4226_ (.A1(_0896_),
    .A2(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4227_ (.A1(_0892_),
    .A2(_0901_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4228_ (.A1(_0892_),
    .A2(_0901_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4229_ (.A1(_0902_),
    .A2(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4230_ (.I(_0843_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4231_ (.A1(_0841_),
    .A2(_0850_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4232_ (.A1(_0841_),
    .A2(_0850_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4233_ (.A1(_0905_),
    .A2(_0906_),
    .B(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4234_ (.A1(_0666_),
    .A2(_0849_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4235_ (.A1(_0655_),
    .A2(_0665_),
    .A3(\mod.Arithmetic.CN.I_in[64] ),
    .A4(_0849_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4236_ (.A1(_0845_),
    .A2(_0909_),
    .B(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4237_ (.A1(_0670_),
    .A2(_0848_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4238_ (.A1(_0671_),
    .A2(_0848_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4239_ (.A1(_0846_),
    .A2(_0912_),
    .A3(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4240_ (.A1(_0641_),
    .A2(\mod.Arithmetic.CN.I_in[66] ),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4241_ (.A1(_0648_),
    .A2(\mod.Arithmetic.ACTI.x[1] ),
    .A3(_0669_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4242_ (.A1(_0647_),
    .A2(\mod.Arithmetic.ACTI.x[2] ),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4243_ (.A1(_0846_),
    .A2(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4244_ (.A1(_0916_),
    .A2(_0918_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4245_ (.A1(_0912_),
    .A2(_0915_),
    .A3(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4246_ (.A1(_0914_),
    .A2(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4247_ (.I(\mod.Arithmetic.CN.I_in[58] ),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4248_ (.I(_0922_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4249_ (.A1(_0655_),
    .A2(\mod.Arithmetic.CN.I_in[57] ),
    .A3(_0663_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4250_ (.A1(_0620_),
    .A2(_0922_),
    .A3(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4251_ (.A1(_0923_),
    .A2(_0924_),
    .B(_0925_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4252_ (.A1(_0911_),
    .A2(_0921_),
    .A3(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4253_ (.I(\mod.Arithmetic.CN.I_in[50] ),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4254_ (.I(_0928_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4255_ (.I(\mod.Arithmetic.CN.I_in[49] ),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4256_ (.A1(_0828_),
    .A2(_0930_),
    .A3(_0660_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4257_ (.A1(_0828_),
    .A2(_0929_),
    .A3(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4258_ (.A1(_0929_),
    .A2(_0931_),
    .B(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4259_ (.A1(_0908_),
    .A2(_0927_),
    .A3(_0933_),
    .Z(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4260_ (.A1(_0891_),
    .A2(_0904_),
    .A3(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4261_ (.A1(_0868_),
    .A2(_0888_),
    .A3(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4262_ (.A1(_0867_),
    .A2(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4263_ (.A1(_0864_),
    .A2(_0937_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4264_ (.A1(_0863_),
    .A2(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4265_ (.I0(_0774_),
    .I1(_0779_),
    .S(_0800_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4266_ (.A1(_0774_),
    .A2(_0857_),
    .B1(_0859_),
    .B2(_0940_),
    .C(_0627_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4267_ (.A1(_0629_),
    .A2(_0939_),
    .B(_0941_),
    .ZN(\mod.P3.Res[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4268_ (.A1(_0863_),
    .A2(_0938_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4269_ (.I(_0864_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4270_ (.A1(_0867_),
    .A2(_0936_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4271_ (.A1(_0943_),
    .A2(_0937_),
    .B(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4272_ (.A1(_0869_),
    .A2(_0887_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4273_ (.A1(_0868_),
    .A2(_0888_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4274_ (.A1(_0946_),
    .A2(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4275_ (.A1(_0868_),
    .A2(_0888_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4276_ (.A1(_0904_),
    .A2(_0934_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4277_ (.A1(_0947_),
    .A2(_0949_),
    .A3(_0935_),
    .B1(_0950_),
    .B2(_0891_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4278_ (.A1(_0883_),
    .A2(_0886_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4279_ (.A1(_0693_),
    .A2(_0810_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4280_ (.A1(_0873_),
    .A2(_0650_),
    .A3(_0813_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4281_ (.A1(_0879_),
    .A2(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4282_ (.A1(_0667_),
    .A2(\mod.Arithmetic.CN.I_in[19] ),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4283_ (.A1(_0877_),
    .A2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4284_ (.I(\mod.Arithmetic.CN.I_in[27] ),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4285_ (.I(_0958_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4286_ (.A1(_0959_),
    .A2(_0812_),
    .A3(_0875_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4287_ (.A1(_0648_),
    .A2(_0959_),
    .B1(_0812_),
    .B2(_0875_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4288_ (.A1(_0957_),
    .A2(_0960_),
    .A3(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4289_ (.A1(_0960_),
    .A2(_0961_),
    .B(_0957_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4290_ (.A1(_0962_),
    .A2(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4291_ (.A1(_0953_),
    .A2(_0955_),
    .A3(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4292_ (.A1(_0872_),
    .A2(_0880_),
    .A3(_0881_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4293_ (.A1(_0880_),
    .A2(_0881_),
    .B(_0872_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4294_ (.A1(_0870_),
    .A2(_0966_),
    .A3(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4295_ (.A1(_0966_),
    .A2(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4296_ (.A1(_0965_),
    .A2(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4297_ (.A1(_0618_),
    .A2(\mod.Arithmetic.CN.I_in[11] ),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4298_ (.I(_0971_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4299_ (.A1(_0722_),
    .A2(_0820_),
    .B1(_0884_),
    .B2(_0715_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4300_ (.A1(_0972_),
    .A2(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4301_ (.A1(_0902_),
    .A2(_0970_),
    .A3(_0974_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4302_ (.A1(_0952_),
    .A2(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4303_ (.A1(_0927_),
    .A2(_0933_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4304_ (.A1(_0902_),
    .A2(_0903_),
    .A3(_0934_),
    .B1(_0977_),
    .B2(_0908_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4305_ (.A1(_0896_),
    .A2(_0900_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4306_ (.A1(_0644_),
    .A2(\mod.Arithmetic.CN.I_in[35] ),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4307_ (.A1(_0894_),
    .A2(_0832_),
    .B1(_0893_),
    .B2(\mod.Arithmetic.CN.I_in[33] ),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4308_ (.A1(_0980_),
    .A2(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4309_ (.A1(_0634_),
    .A2(\mod.Arithmetic.CN.I_in[43] ),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4310_ (.I(_0983_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4311_ (.A1(_0898_),
    .A2(_0837_),
    .B1(_0897_),
    .B2(\mod.Arithmetic.CN.I_in[41] ),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4312_ (.A1(_0984_),
    .A2(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4313_ (.A1(_0982_),
    .A2(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4314_ (.A1(_0979_),
    .A2(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4315_ (.A1(_0979_),
    .A2(_0987_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4316_ (.A1(_0988_),
    .A2(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4317_ (.A1(_0921_),
    .A2(_0926_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4318_ (.A1(_0911_),
    .A2(_0991_),
    .B1(_0927_),
    .B2(_0933_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4319_ (.A1(_0929_),
    .A2(_0660_),
    .A3(_0842_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4320_ (.A1(_0922_),
    .A2(_0663_),
    .A3(_0844_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4321_ (.A1(_0658_),
    .A2(_0928_),
    .A3(\mod.Arithmetic.CN.I_in[51] ),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4322_ (.A1(_0658_),
    .A2(\mod.Arithmetic.CN.I_in[50] ),
    .A3(_0842_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4323_ (.A1(_0649_),
    .A2(\mod.Arithmetic.CN.I_in[51] ),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4324_ (.A1(_0930_),
    .A2(_0995_),
    .B1(_0996_),
    .B2(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4325_ (.A1(_0994_),
    .A2(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4326_ (.A1(_0993_),
    .A2(_0999_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4327_ (.A1(_0993_),
    .A2(_0999_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4328_ (.A1(_1000_),
    .A2(_1001_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4329_ (.A1(_0914_),
    .A2(_0920_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4330_ (.A1(_0921_),
    .A2(_0926_),
    .B(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4331_ (.A1(_0912_),
    .A2(_0919_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4332_ (.A1(_0671_),
    .A2(_0848_),
    .A3(_0919_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4333_ (.A1(_0915_),
    .A2(_1005_),
    .B(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4334_ (.A1(_0646_),
    .A2(\mod.Arithmetic.CN.I_in[67] ),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4335_ (.A1(\mod.Arithmetic.CN.I_in[64] ),
    .A2(_0918_),
    .B(\mod.Arithmetic.ACTI.x[1] ),
    .C(_0634_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4336_ (.A1(_0633_),
    .A2(\mod.Arithmetic.ACTI.x[2] ),
    .A3(_0846_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4337_ (.A1(_0615_),
    .A2(\mod.Arithmetic.ACTI.x[3] ),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4338_ (.A1(_0915_),
    .A2(_1011_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4339_ (.A1(_1010_),
    .A2(_1012_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4340_ (.A1(_1009_),
    .A2(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4341_ (.A1(_1008_),
    .A2(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4342_ (.A1(_1007_),
    .A2(_1015_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4343_ (.I(\mod.Arithmetic.CN.I_in[59] ),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4344_ (.I(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4345_ (.A1(_0649_),
    .A2(_1017_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4346_ (.A1(_0817_),
    .A2(_0923_),
    .A3(_0844_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4347_ (.I0(_1018_),
    .I1(_1019_),
    .S(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4348_ (.A1(_1004_),
    .A2(_1016_),
    .A3(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4349_ (.A1(_0992_),
    .A2(_1002_),
    .A3(_1022_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4350_ (.A1(_0978_),
    .A2(_0990_),
    .A3(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4351_ (.A1(_0951_),
    .A2(_0976_),
    .A3(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4352_ (.A1(_0948_),
    .A2(_1025_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4353_ (.A1(_0945_),
    .A2(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4354_ (.A1(_0942_),
    .A2(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4355_ (.I0(_0781_),
    .I1(_0780_),
    .S(_0800_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4356_ (.A1(_0781_),
    .A2(_0857_),
    .B1(_0858_),
    .B2(_1029_),
    .C(_0627_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4357_ (.A1(_0629_),
    .A2(_1028_),
    .B(_1030_),
    .ZN(\mod.P3.Res[3] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4358_ (.I(_0627_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4359_ (.A1(_0787_),
    .A2(_0805_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4360_ (.A1(_0786_),
    .A2(_0801_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4361_ (.A1(_0787_),
    .A2(_0856_),
    .B1(_0858_),
    .B2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4362_ (.A1(_0945_),
    .A2(_1026_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4363_ (.A1(_0863_),
    .A2(_0938_),
    .A3(_1027_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4364_ (.A1(_0976_),
    .A2(_1024_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4365_ (.A1(_0948_),
    .A2(_1025_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4366_ (.A1(_0951_),
    .A2(_1037_),
    .B(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4367_ (.A1(_0970_),
    .A2(_0974_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4368_ (.A1(_0902_),
    .A2(_1040_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4369_ (.A1(_0952_),
    .A2(_0975_),
    .B(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4370_ (.A1(_0990_),
    .A2(_1023_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4371_ (.A1(_0978_),
    .A2(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4372_ (.A1(_0976_),
    .A2(_1024_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4373_ (.A1(_1044_),
    .A2(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4374_ (.A1(_0970_),
    .A2(_0974_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4375_ (.A1(_0968_),
    .A2(_0965_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4376_ (.A1(_0966_),
    .A2(_0965_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4377_ (.A1(_0962_),
    .A2(_0963_),
    .B(_0879_),
    .C(_0954_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4378_ (.A1(_0880_),
    .A2(_0954_),
    .B(_0962_),
    .C(_0963_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4379_ (.A1(_0693_),
    .A2(_0810_),
    .A3(_1050_),
    .B(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4380_ (.A1(_0617_),
    .A2(_0686_),
    .A3(_0688_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4381_ (.A1(_0957_),
    .A2(_0960_),
    .A3(_0961_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4382_ (.A1(_0668_),
    .A2(\mod.Arithmetic.CN.I_in[26] ),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4383_ (.A1(_0643_),
    .A2(_0959_),
    .B(_0813_),
    .C(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4384_ (.A1(_1054_),
    .A2(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4385_ (.A1(_0616_),
    .A2(_0697_),
    .A3(\mod.Arithmetic.CN.I_in[19] ),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4386_ (.A1(_0640_),
    .A2(\mod.Arithmetic.CN.I_in[20] ),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4387_ (.A1(_0956_),
    .A2(_1059_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4388_ (.I(_0640_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4389_ (.I(\mod.Arithmetic.CN.I_in[28] ),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4390_ (.I(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4391_ (.A1(_0613_),
    .A2(\mod.Arithmetic.CN.I_in[27] ),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4392_ (.A1(_1061_),
    .A2(_1063_),
    .B1(_1064_),
    .B2(_0873_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4393_ (.A1(_0633_),
    .A2(_0959_),
    .A3(_1062_),
    .A4(_1055_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4394_ (.A1(_1058_),
    .A2(_1060_),
    .A3(_1065_),
    .A4(_1066_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4395_ (.A1(_0956_),
    .A2(_1059_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4396_ (.A1(_0647_),
    .A2(_0958_),
    .A3(_1063_),
    .A4(_1055_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4397_ (.A1(_0639_),
    .A2(\mod.Arithmetic.CN.I_in[28] ),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4398_ (.A1(\mod.Arithmetic.CN.I_in[26] ),
    .A2(_1064_),
    .B(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4399_ (.A1(_1068_),
    .A2(_1069_),
    .A3(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4400_ (.A1(_1067_),
    .A2(_1072_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4401_ (.A1(_1053_),
    .A2(_1057_),
    .A3(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4402_ (.A1(_1052_),
    .A2(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4403_ (.A1(_0894_),
    .A2(_0832_),
    .A3(_0980_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4404_ (.A1(_1049_),
    .A2(_1075_),
    .A3(_1076_),
    .Z(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4405_ (.A1(_0620_),
    .A2(_0730_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4406_ (.A1(_0620_),
    .A2(_0728_),
    .A3(_0721_),
    .A4(\mod.Arithmetic.CN.I_in[9] ),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4407_ (.A1(_0721_),
    .A2(_0972_),
    .B(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4408_ (.A1(_0722_),
    .A2(_0820_),
    .A3(_0972_),
    .B(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4409_ (.A1(_1078_),
    .A2(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4410_ (.A1(_1048_),
    .A2(_1077_),
    .A3(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4411_ (.A1(_0988_),
    .A2(_1083_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4412_ (.A1(_1002_),
    .A2(_1022_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4413_ (.A1(_1002_),
    .A2(_1022_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _4414_ (.A1(_0992_),
    .A2(_1085_),
    .A3(_1086_),
    .B1(_1023_),
    .B2(_0988_),
    .B3(_0989_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4415_ (.I(_0986_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4416_ (.A1(_0982_),
    .A2(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4417_ (.I(\mod.Arithmetic.CN.I_in[36] ),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4418_ (.A1(_0619_),
    .A2(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4419_ (.A1(_0894_),
    .A2(_0980_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4420_ (.A1(_0834_),
    .A2(\mod.Arithmetic.CN.I_in[35] ),
    .B(_0830_),
    .C(_0893_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4421_ (.A1(_1092_),
    .A2(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4422_ (.A1(_1091_),
    .A2(_1094_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4423_ (.A1(_0664_),
    .A2(\mod.Arithmetic.CN.I_in[44] ),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4424_ (.A1(_0898_),
    .A2(_0984_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4425_ (.A1(_0834_),
    .A2(\mod.Arithmetic.CN.I_in[41] ),
    .A3(_0898_),
    .A4(_0984_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4426_ (.A1(_0837_),
    .A2(_1097_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4427_ (.A1(_1097_),
    .A2(_1098_),
    .B(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4428_ (.A1(_1096_),
    .A2(_1100_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4429_ (.A1(_1095_),
    .A2(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4430_ (.A1(_1089_),
    .A2(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4431_ (.A1(_0828_),
    .A2(_1018_),
    .A3(_1020_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4432_ (.A1(_1018_),
    .A2(_1020_),
    .B(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4433_ (.A1(_1004_),
    .A2(_1016_),
    .A3(_1105_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4434_ (.A1(_1016_),
    .A2(_1021_),
    .Z(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4435_ (.A1(_1000_),
    .A2(_1001_),
    .A3(_1106_),
    .B1(_1107_),
    .B2(_1004_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4436_ (.A1(_0930_),
    .A2(_0995_),
    .B1(_0996_),
    .B2(_0997_),
    .C(_0994_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4437_ (.A1(_0993_),
    .A2(_0999_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4438_ (.A1(_1109_),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4439_ (.A1(_0644_),
    .A2(\mod.Arithmetic.CN.I_in[57] ),
    .A3(_0922_),
    .A4(_1019_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4440_ (.A1(\mod.Arithmetic.CN.I_in[52] ),
    .A2(_0997_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(_0642_),
    .A2(\mod.Arithmetic.CN.I_in[51] ),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4442_ (.A1(\mod.Arithmetic.CN.I_in[50] ),
    .A2(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4443_ (.A1(_0632_),
    .A2(\mod.Arithmetic.CN.I_in[52] ),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4444_ (.A1(_0928_),
    .A2(_1113_),
    .B1(_1115_),
    .B2(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4445_ (.A1(_1112_),
    .A2(_1117_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4446_ (.A1(_0619_),
    .A2(_0930_),
    .A3(_0928_),
    .A4(_1114_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4447_ (.A1(_1118_),
    .A2(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4448_ (.A1(_1111_),
    .A2(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4449_ (.A1(_1007_),
    .A2(_1015_),
    .B1(_1016_),
    .B2(_1105_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4450_ (.A1(_1009_),
    .A2(_1013_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4451_ (.A1(_1008_),
    .A2(_1014_),
    .B(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4452_ (.A1(_0667_),
    .A2(\mod.Arithmetic.CN.I_in[68] ),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4453_ (.A1(\mod.Arithmetic.CN.I_in[65] ),
    .A2(_1012_),
    .B(_0643_),
    .C(\mod.Arithmetic.ACTI.x[2] ),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4454_ (.A1(_0642_),
    .A2(\mod.Arithmetic.ACTI.x[3] ),
    .A3(_0915_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4455_ (.A1(_0614_),
    .A2(\mod.Arithmetic.ACTI.x[4] ),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4456_ (.A1(_1008_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4457_ (.A1(_1127_),
    .A2(_1129_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4458_ (.A1(_1126_),
    .A2(_1130_),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4459_ (.A1(_1125_),
    .A2(_1131_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4460_ (.A1(_1124_),
    .A2(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4461_ (.I(\mod.Arithmetic.CN.I_in[60] ),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4462_ (.A1(_0661_),
    .A2(_1017_),
    .A3(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4463_ (.A1(_0616_),
    .A2(\mod.Arithmetic.CN.I_in[60] ),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4464_ (.A1(_0923_),
    .A2(_1019_),
    .B(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4465_ (.A1(_0923_),
    .A2(_1135_),
    .B(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4466_ (.A1(_1133_),
    .A2(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4467_ (.A1(_1121_),
    .A2(_1122_),
    .A3(_1139_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4468_ (.A1(_1103_),
    .A2(_1108_),
    .A3(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4469_ (.A1(_1087_),
    .A2(_1141_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4470_ (.A1(_1047_),
    .A2(_1084_),
    .A3(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4471_ (.A1(_1042_),
    .A2(_1046_),
    .A3(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4472_ (.A1(_1039_),
    .A2(_1144_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4473_ (.A1(_1035_),
    .A2(_1036_),
    .A3(_1145_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4474_ (.A1(_1035_),
    .A2(_1036_),
    .B(_1145_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4475_ (.A1(_1031_),
    .A2(_1146_),
    .A3(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4476_ (.A1(_1031_),
    .A2(_1032_),
    .A3(_1034_),
    .B(_1148_),
    .ZN(\mod.P3.Res[4] ));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4477_ (.A1(_0731_),
    .A2(_0722_),
    .A3(_0820_),
    .A4(_0972_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4478_ (.A1(_1044_),
    .A2(_1045_),
    .A3(_1143_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4479_ (.A1(_1044_),
    .A2(_1045_),
    .B(_1143_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4480_ (.A1(_1042_),
    .A2(_1150_),
    .B(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4481_ (.A1(_1047_),
    .A2(_1084_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4482_ (.A1(_0988_),
    .A2(_1083_),
    .B(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4483_ (.A1(_1047_),
    .A2(_1084_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4484_ (.A1(_1087_),
    .A2(_1141_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4485_ (.A1(_1087_),
    .A2(_1141_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4486_ (.A1(_1153_),
    .A2(_1155_),
    .A3(_1156_),
    .B(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4487_ (.A1(_1089_),
    .A2(_1102_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4488_ (.A1(_1048_),
    .A2(_1077_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4489_ (.A1(_1048_),
    .A2(_1077_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4490_ (.A1(_1160_),
    .A2(_1082_),
    .B(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4491_ (.A1(_1075_),
    .A2(_1076_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4492_ (.A1(_1075_),
    .A2(_1076_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4493_ (.A1(_1049_),
    .A2(_1163_),
    .B(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4494_ (.A1(_1052_),
    .A2(_1074_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4495_ (.A1(_1067_),
    .A2(_1072_),
    .B(_1054_),
    .C(_1056_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4496_ (.A1(_1054_),
    .A2(_1056_),
    .B(_1067_),
    .C(_1072_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4497_ (.A1(_1053_),
    .A2(_1167_),
    .B(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4498_ (.A1(_1069_),
    .A2(_1071_),
    .B(_1068_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4499_ (.A1(_1055_),
    .A2(_1064_),
    .A3(_1070_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4500_ (.A1(_1170_),
    .A2(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4501_ (.A1(_0684_),
    .A2(\mod.Arithmetic.CN.I_in[20] ),
    .B(_0613_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4502_ (.A1(_0639_),
    .A2(\mod.Arithmetic.CN.I_in[21] ),
    .A3(\mod.Arithmetic.CN.I_in[20] ),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4503_ (.A1(_1173_),
    .A2(_1174_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4504_ (.A1(_0613_),
    .A2(_1062_),
    .A3(\mod.Arithmetic.CN.I_in[29] ),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4505_ (.A1(_0958_),
    .A2(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4506_ (.I(\mod.Arithmetic.CN.I_in[29] ),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4507_ (.A1(_0646_),
    .A2(_1178_),
    .B1(_1064_),
    .B2(_1070_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4508_ (.A1(_1175_),
    .A2(_1177_),
    .A3(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4509_ (.A1(_1177_),
    .A2(_1179_),
    .B(_1175_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4510_ (.A1(_1180_),
    .A2(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4511_ (.A1(_1058_),
    .A2(_1172_),
    .A3(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4512_ (.A1(_1169_),
    .A2(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4513_ (.I(_1090_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4514_ (.A1(_1185_),
    .A2(_1093_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4515_ (.A1(_1166_),
    .A2(_1184_),
    .A3(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4516_ (.A1(_0621_),
    .A2(_0737_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4517_ (.I(\mod.Arithmetic.CN.I_in[12] ),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4518_ (.I(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4519_ (.A1(_0730_),
    .A2(_0713_),
    .A3(_0971_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4520_ (.A1(\mod.Arithmetic.CN.I_in[11] ),
    .A2(_1078_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4521_ (.A1(_1190_),
    .A2(_1079_),
    .B1(_1191_),
    .B2(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4522_ (.A1(_1188_),
    .A2(_1193_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4523_ (.I(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4524_ (.A1(_1165_),
    .A2(_1187_),
    .A3(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4525_ (.A1(_1159_),
    .A2(_1162_),
    .A3(_1196_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4526_ (.I(_1103_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4527_ (.A1(_1108_),
    .A2(_1140_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4528_ (.A1(_1108_),
    .A2(_1140_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4529_ (.A1(_1198_),
    .A2(_1199_),
    .B(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4530_ (.I(\mod.Arithmetic.CN.I_in[44] ),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4531_ (.I(_1202_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4532_ (.I(_1101_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4533_ (.A1(_1203_),
    .A2(_1099_),
    .B1(_1204_),
    .B2(_1095_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4534_ (.A1(_1203_),
    .A2(_1098_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4535_ (.I(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4536_ (.I(\mod.Arithmetic.CN.I_in[45] ),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4537_ (.A1(_0659_),
    .A2(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4538_ (.A1(_0664_),
    .A2(\mod.Arithmetic.CN.I_in[44] ),
    .B(_0897_),
    .C(_0983_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4539_ (.A1(\mod.Arithmetic.CN.I_in[43] ),
    .A2(_1096_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4540_ (.A1(_1210_),
    .A2(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4541_ (.A1(_1209_),
    .A2(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4542_ (.A1(_0636_),
    .A2(\mod.Arithmetic.CN.I_in[37] ),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4543_ (.A1(_0635_),
    .A2(\mod.Arithmetic.CN.I_in[36] ),
    .B(_0893_),
    .C(_0980_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4544_ (.A1(\mod.Arithmetic.CN.I_in[35] ),
    .A2(_1091_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4545_ (.A1(_1215_),
    .A2(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4546_ (.A1(_1214_),
    .A2(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4547_ (.A1(_1207_),
    .A2(_1213_),
    .A3(_1218_),
    .Z(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4548_ (.A1(_1205_),
    .A2(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4549_ (.A1(_1122_),
    .A2(_1139_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4550_ (.A1(_1122_),
    .A2(_1139_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4551_ (.A1(_1121_),
    .A2(_1221_),
    .B(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4552_ (.A1(_0929_),
    .A2(_1113_),
    .B1(_1115_),
    .B2(_1116_),
    .C(_1112_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4553_ (.A1(_1118_),
    .A2(_1119_),
    .B(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(\mod.Arithmetic.CN.I_in[52] ),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4555_ (.A1(_1226_),
    .A2(_0995_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4556_ (.A1(_0643_),
    .A2(\mod.Arithmetic.CN.I_in[58] ),
    .A3(\mod.Arithmetic.CN.I_in[59] ),
    .A4(_1136_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4557_ (.A1(_0633_),
    .A2(\mod.Arithmetic.CN.I_in[53] ),
    .B1(_1114_),
    .B2(_1116_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4558_ (.A1(\mod.Arithmetic.CN.I_in[53] ),
    .A2(_1114_),
    .A3(_1116_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4559_ (.A1(_1229_),
    .A2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4560_ (.A1(_1228_),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4561_ (.A1(_1227_),
    .A2(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4562_ (.A1(_1225_),
    .A2(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4563_ (.A1(_1111_),
    .A2(_1120_),
    .A3(_1234_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4564_ (.A1(_1111_),
    .A2(_1120_),
    .B(_1234_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4565_ (.A1(_1235_),
    .A2(_1236_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4566_ (.A1(_1124_),
    .A2(_1132_),
    .B1(_1133_),
    .B2(_1138_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4567_ (.A1(_0664_),
    .A2(\mod.Arithmetic.CN.I_in[68] ),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4568_ (.A1(_1126_),
    .A2(_1130_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4569_ (.A1(_1239_),
    .A2(_1131_),
    .B(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4570_ (.A1(_0667_),
    .A2(\mod.Arithmetic.CN.I_in[69] ),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4571_ (.A1(\mod.Arithmetic.CN.I_in[66] ),
    .A2(_1129_),
    .B(_0648_),
    .C(_0781_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4572_ (.A1(\mod.Arithmetic.CN.I_in[67] ),
    .A2(_1128_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4573_ (.A1(_0640_),
    .A2(\mod.Arithmetic.ACTI.x[5] ),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4574_ (.A1(_1125_),
    .A2(_1245_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4575_ (.A1(_1244_),
    .A2(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4576_ (.A1(_1243_),
    .A2(_1247_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4577_ (.A1(_1242_),
    .A2(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4578_ (.A1(_1241_),
    .A2(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4579_ (.I(\mod.Arithmetic.CN.I_in[61] ),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4580_ (.I(_1061_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4581_ (.A1(_1252_),
    .A2(_1251_),
    .B1(_1136_),
    .B2(_1017_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4582_ (.A1(_1018_),
    .A2(_1251_),
    .A3(_1136_),
    .B(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4583_ (.A1(_1250_),
    .A2(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4584_ (.A1(_1238_),
    .A2(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4585_ (.A1(_1237_),
    .A2(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4586_ (.A1(_1220_),
    .A2(_1223_),
    .A3(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4587_ (.A1(_1197_),
    .A2(_1201_),
    .A3(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4588_ (.A1(_1154_),
    .A2(_1158_),
    .A3(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4589_ (.A1(_1149_),
    .A2(_1152_),
    .A3(_1260_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4590_ (.A1(_1039_),
    .A2(_1144_),
    .B(_1147_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4591_ (.A1(_1261_),
    .A2(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4592_ (.A1(_0791_),
    .A2(_0801_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4593_ (.A1(_0792_),
    .A2(_0805_),
    .B(_0859_),
    .C(_1264_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4594_ (.A1(_0792_),
    .A2(_0857_),
    .B(_0628_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4595_ (.A1(_1031_),
    .A2(_1263_),
    .B1(_1265_),
    .B2(_1266_),
    .ZN(\mod.P3.Res[5] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4596_ (.A1(_0805_),
    .A2(_0859_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4597_ (.A1(\mod.P2.Rout_reg[0] ),
    .A2(_0678_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4598_ (.A1(\mod.Arithmetic.ACTI.x[6] ),
    .A2(_1268_),
    .A3(_0802_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4599_ (.A1(_1261_),
    .A2(_1262_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4600_ (.A1(_1152_),
    .A2(_1260_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4601_ (.A1(_1152_),
    .A2(_1260_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4602_ (.A1(_1149_),
    .A2(_1271_),
    .B(_1272_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4603_ (.A1(_0625_),
    .A2(_0738_),
    .B(_1190_),
    .C(_1079_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4604_ (.A1(_1158_),
    .A2(_1259_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4605_ (.A1(_1158_),
    .A2(_1259_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4606_ (.A1(_1154_),
    .A2(_1275_),
    .B(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4607_ (.A1(_1159_),
    .A2(_1196_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4608_ (.A1(_1162_),
    .A2(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4609_ (.A1(_1159_),
    .A2(_1196_),
    .B(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4610_ (.A1(_1201_),
    .A2(_1258_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4611_ (.A1(_1201_),
    .A2(_1258_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4612_ (.A1(_1197_),
    .A2(_1281_),
    .B(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4613_ (.A1(_1165_),
    .A2(_1187_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4614_ (.A1(_1165_),
    .A2(_1187_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4615_ (.A1(_1284_),
    .A2(_1195_),
    .B(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4616_ (.A1(_1205_),
    .A2(_1219_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4617_ (.I(\mod.Arithmetic.CN.I_in[13] ),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4618_ (.I(\mod.Arithmetic.CN.I_in[14] ),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4619_ (.A1(_1288_),
    .A2(_0730_),
    .B(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4620_ (.A1(_0743_),
    .A2(\mod.Arithmetic.CN.I_in[13] ),
    .A3(_1190_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4621_ (.A1(_0834_),
    .A2(_1290_),
    .A3(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4622_ (.A1(_0737_),
    .A2(_1191_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4623_ (.A1(_1292_),
    .A2(_1293_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4624_ (.A1(\mod.Arithmetic.CN.I_in[13] ),
    .A2(_1189_),
    .A3(_0971_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4625_ (.I0(_1292_),
    .I1(_0743_),
    .S(_1295_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4626_ (.A1(_1293_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4627_ (.A1(_1294_),
    .A2(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4628_ (.A1(_1185_),
    .A2(_1093_),
    .B(_1184_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4629_ (.A1(_1185_),
    .A2(_1093_),
    .A3(_1184_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4630_ (.A1(_1166_),
    .A2(_1299_),
    .B(_1300_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4631_ (.A1(_1169_),
    .A2(_1183_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4632_ (.I(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4633_ (.A1(\mod.Arithmetic.CN.I_in[37] ),
    .A2(_1215_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4634_ (.A1(_1180_),
    .A2(_1181_),
    .B(_1170_),
    .C(_1171_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4635_ (.A1(_1170_),
    .A2(_1171_),
    .B(_1180_),
    .C(_1181_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4636_ (.A1(_1058_),
    .A2(_1305_),
    .B(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4637_ (.I(_1178_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4638_ (.A1(_0647_),
    .A2(_0958_),
    .A3(_1062_),
    .A4(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4639_ (.A1(_1180_),
    .A2(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4640_ (.A1(_0614_),
    .A2(\mod.Arithmetic.CN.I_in[22] ),
    .A3(_0684_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4641_ (.A1(_0701_),
    .A2(_0685_),
    .B(_1061_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4642_ (.A1(_1311_),
    .A2(_1312_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4643_ (.A1(_1063_),
    .A2(_1178_),
    .A3(\mod.Arithmetic.CN.I_in[30] ),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4644_ (.I(\mod.Arithmetic.CN.I_in[30] ),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4645_ (.A1(_1063_),
    .A2(_1178_),
    .B(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4646_ (.A1(_1061_),
    .A2(_1314_),
    .A3(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4647_ (.A1(_1313_),
    .A2(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4648_ (.A1(_1174_),
    .A2(_1310_),
    .A3(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4649_ (.A1(_1307_),
    .A2(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4650_ (.A1(_1304_),
    .A2(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4651_ (.A1(_1303_),
    .A2(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4652_ (.A1(_1298_),
    .A2(_1301_),
    .A3(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4653_ (.A1(_1287_),
    .A2(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4654_ (.A1(_1286_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4655_ (.A1(_1223_),
    .A2(_1257_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4656_ (.A1(_1223_),
    .A2(_1257_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4657_ (.A1(_1220_),
    .A2(_1326_),
    .B(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4658_ (.A1(_1206_),
    .A2(_1213_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4659_ (.A1(_1209_),
    .A2(_1207_),
    .B1(_1329_),
    .B2(_1218_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4660_ (.I(\mod.Arithmetic.CN.I_in[37] ),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4661_ (.A1(_0659_),
    .A2(\mod.Arithmetic.CN.I_in[35] ),
    .A3(_1090_),
    .A4(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4662_ (.A1(_1090_),
    .A2(_1331_),
    .B(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4663_ (.A1(\mod.Arithmetic.CN.I_in[38] ),
    .A2(_1333_),
    .B(_1252_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4664_ (.A1(\mod.Arithmetic.CN.I_in[38] ),
    .A2(_1333_),
    .B(_1334_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4665_ (.A1(_1202_),
    .A2(\mod.Arithmetic.CN.I_in[45] ),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4666_ (.A1(\mod.Arithmetic.CN.I_in[46] ),
    .A2(_1336_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4667_ (.A1(_1252_),
    .A2(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4668_ (.A1(_1203_),
    .A2(\mod.Arithmetic.CN.I_in[45] ),
    .A3(_0984_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4669_ (.A1(\mod.Arithmetic.CN.I_in[46] ),
    .A2(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4670_ (.A1(_1339_),
    .A2(_1338_),
    .B(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4671_ (.A1(_1208_),
    .A2(_1210_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4672_ (.I0(_1338_),
    .I1(_1341_),
    .S(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4673_ (.A1(_1335_),
    .A2(_1343_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4674_ (.A1(_1235_),
    .A2(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4675_ (.A1(_1330_),
    .A2(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4676_ (.I(_1346_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4677_ (.A1(_1238_),
    .A2(_1255_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4678_ (.A1(_1237_),
    .A2(_1256_),
    .B(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4679_ (.A1(_1225_),
    .A2(_1233_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4680_ (.A1(_1228_),
    .A2(_1231_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4681_ (.A1(_1226_),
    .A2(_0995_),
    .A3(_1232_),
    .B(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4682_ (.A1(\mod.Arithmetic.CN.I_in[61] ),
    .A2(_1135_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4683_ (.I(\mod.Arithmetic.CN.I_in[53] ),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4684_ (.A1(\mod.Arithmetic.CN.I_in[52] ),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4685_ (.A1(\mod.Arithmetic.CN.I_in[54] ),
    .A2(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4686_ (.A1(_0618_),
    .A2(_1356_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4687_ (.A1(_1353_),
    .A2(_1356_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4688_ (.A1(_1353_),
    .A2(_1357_),
    .B(_1358_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4689_ (.A1(_1226_),
    .A2(_1354_),
    .A3(_0997_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4690_ (.A1(_1359_),
    .A2(_1360_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4691_ (.A1(_1352_),
    .A2(_1361_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4692_ (.A1(_1350_),
    .A2(_1362_),
    .Z(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4693_ (.A1(_1241_),
    .A2(_1249_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4694_ (.A1(_1250_),
    .A2(_1254_),
    .B(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4695_ (.I(\mod.Arithmetic.CN.I_in[62] ),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4696_ (.A1(_1134_),
    .A2(_1251_),
    .B(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4697_ (.A1(_1134_),
    .A2(_1251_),
    .A3(_1366_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4698_ (.A1(_0636_),
    .A2(_1367_),
    .A3(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4699_ (.A1(_0658_),
    .A2(\mod.Arithmetic.CN.I_in[69] ),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4700_ (.A1(_1243_),
    .A2(_1247_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4701_ (.A1(_1370_),
    .A2(_1248_),
    .B(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4702_ (.A1(_0661_),
    .A2(\mod.Arithmetic.CN.I_in[70] ),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4703_ (.A1(\mod.Arithmetic.CN.I_in[67] ),
    .A2(_1246_),
    .B(_0642_),
    .C(\mod.Arithmetic.ACTI.x[4] ),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4704_ (.A1(_0641_),
    .A2(\mod.Arithmetic.ACTI.x[5] ),
    .A3(_1125_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4705_ (.A1(_0646_),
    .A2(\mod.Arithmetic.ACTI.x[6] ),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4706_ (.A1(_1242_),
    .A2(_1376_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4707_ (.A1(_1375_),
    .A2(_1377_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4708_ (.A1(_1374_),
    .A2(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4709_ (.A1(_1373_),
    .A2(_1379_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4710_ (.A1(_1372_),
    .A2(_1380_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4711_ (.A1(_1369_),
    .A2(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4712_ (.A1(_1365_),
    .A2(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4713_ (.A1(_1363_),
    .A2(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4714_ (.A1(_1349_),
    .A2(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4715_ (.A1(_1347_),
    .A2(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4716_ (.A1(_1325_),
    .A2(_1328_),
    .A3(_1386_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4717_ (.A1(_1280_),
    .A2(_1283_),
    .A3(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4718_ (.A1(_1277_),
    .A2(_1388_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4719_ (.A1(_1274_),
    .A2(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4720_ (.A1(_1273_),
    .A2(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4721_ (.A1(_1270_),
    .A2(_1391_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4722_ (.A1(_1270_),
    .A2(_1391_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4723_ (.A1(_1031_),
    .A2(_1392_),
    .A3(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4724_ (.A1(_0795_),
    .A2(_1267_),
    .B(_1269_),
    .C(_1394_),
    .ZN(\mod.P3.Res[6] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4725_ (.A1(_1273_),
    .A2(_1390_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4726_ (.A1(_1277_),
    .A2(_1388_),
    .B1(_1389_),
    .B2(_1274_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4727_ (.A1(_1283_),
    .A2(_1387_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4728_ (.A1(_1283_),
    .A2(_1387_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4729_ (.A1(_1280_),
    .A2(_1397_),
    .B(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4730_ (.I(_1349_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4731_ (.A1(_1347_),
    .A2(_1385_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4732_ (.A1(_1400_),
    .A2(_1384_),
    .B(_1401_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4733_ (.A1(\mod.Arithmetic.CN.I_in[61] ),
    .A2(_1366_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4734_ (.A1(\mod.Arithmetic.CN.I_in[63] ),
    .A2(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4735_ (.A1(_0625_),
    .A2(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4736_ (.A1(_1294_),
    .A2(_1402_),
    .A3(_1405_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4737_ (.A1(_1350_),
    .A2(_1362_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4738_ (.A1(_1208_),
    .A2(_1210_),
    .A3(_1338_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4739_ (.A1(_1335_),
    .A2(_1343_),
    .B(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4740_ (.A1(_1407_),
    .A2(_1409_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4741_ (.I(_1208_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4742_ (.A1(_1411_),
    .A2(\mod.Arithmetic.CN.I_in[46] ),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4743_ (.A1(\mod.Arithmetic.CN.I_in[47] ),
    .A2(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4744_ (.A1(_0622_),
    .A2(_1413_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4745_ (.A1(_0622_),
    .A2(\mod.Arithmetic.CN.I_in[71] ),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4746_ (.A1(\mod.Arithmetic.CN.I_in[69] ),
    .A2(_1376_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4747_ (.I0(_1373_),
    .I1(\mod.Arithmetic.CN.I_in[70] ),
    .S(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4748_ (.A1(_1414_),
    .A2(_1415_),
    .A3(_1417_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4749_ (.A1(_0623_),
    .A2(\mod.Arithmetic.CN.I_in[70] ),
    .A3(_1379_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4750_ (.A1(_1374_),
    .A2(_1378_),
    .B(_1419_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4751_ (.A1(_1203_),
    .A2(\mod.Arithmetic.CN.I_in[46] ),
    .A3(_1209_),
    .B(_1340_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4752_ (.I(_0622_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4753_ (.I(\mod.Arithmetic.CN.I_in[38] ),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4754_ (.A1(_1185_),
    .A2(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4755_ (.A1(\mod.Arithmetic.CN.I_in[37] ),
    .A2(_1423_),
    .B1(_1214_),
    .B2(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4756_ (.A1(\mod.Arithmetic.CN.I_in[39] ),
    .A2(_1425_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4757_ (.A1(_1422_),
    .A2(_1426_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4758_ (.A1(_1421_),
    .A2(_1427_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4759_ (.A1(_1418_),
    .A2(_1420_),
    .A3(_1428_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4760_ (.A1(_1287_),
    .A2(_1323_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4761_ (.A1(_1286_),
    .A2(_1324_),
    .B(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4762_ (.A1(_1410_),
    .A2(_1429_),
    .A3(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4763_ (.A1(_1252_),
    .A2(_1354_),
    .A3(\mod.Arithmetic.CN.I_in[54] ),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4764_ (.A1(_1352_),
    .A2(_1361_),
    .B1(_1433_),
    .B2(_1226_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4765_ (.A1(_1359_),
    .A2(_1360_),
    .B(_1434_),
    .C(_1358_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4766_ (.A1(_1422_),
    .A2(\mod.Arithmetic.ACTI.x[7] ),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4767_ (.A1(\mod.Arithmetic.CN.I_in[68] ),
    .A2(_1377_),
    .B(_1422_),
    .C(\mod.Arithmetic.ACTI.x[5] ),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4768_ (.I0(\mod.Arithmetic.ACTI.x[7] ),
    .I1(_1436_),
    .S(_1437_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4769_ (.A1(_0624_),
    .A2(_1134_),
    .A3(\mod.Arithmetic.CN.I_in[61] ),
    .A4(_1366_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4770_ (.A1(_0624_),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4771_ (.A1(_1354_),
    .A2(\mod.Arithmetic.CN.I_in[54] ),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4772_ (.A1(\mod.Arithmetic.CN.I_in[55] ),
    .A2(_1441_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4773_ (.I0(_1440_),
    .I1(_1439_),
    .S(_1442_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4774_ (.A1(_1435_),
    .A2(_1438_),
    .A3(_1443_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4775_ (.A1(_1301_),
    .A2(_1322_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4776_ (.A1(_1301_),
    .A2(_1322_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4777_ (.A1(_1298_),
    .A2(_1445_),
    .B(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4778_ (.A1(_1310_),
    .A2(_1318_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4779_ (.A1(_1307_),
    .A2(_1319_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4780_ (.A1(_1310_),
    .A2(_1318_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4781_ (.A1(_1174_),
    .A2(_1448_),
    .B(_1449_),
    .C(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4782_ (.A1(_1447_),
    .A2(_1451_),
    .Z(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4783_ (.A1(_0743_),
    .A2(_1190_),
    .A3(_1188_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4784_ (.A1(_0744_),
    .A2(_1295_),
    .B(_1453_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4785_ (.A1(_1289_),
    .A2(_0737_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4786_ (.A1(\mod.Arithmetic.CN.I_in[15] ),
    .A2(_1455_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4787_ (.A1(_0624_),
    .A2(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4788_ (.A1(_1235_),
    .A2(_1344_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4789_ (.A1(_1330_),
    .A2(_1345_),
    .B(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4790_ (.A1(_1308_),
    .A2(_1315_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4791_ (.A1(\mod.Arithmetic.CN.I_in[23] ),
    .A2(\mod.Arithmetic.CN.I_in[31] ),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4792_ (.A1(_0702_),
    .A2(_1460_),
    .A3(_1461_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4793_ (.A1(_1422_),
    .A2(_1462_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4794_ (.A1(_1423_),
    .A2(_1332_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4795_ (.A1(_1304_),
    .A2(_1320_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4796_ (.A1(_1303_),
    .A2(_1321_),
    .B(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4797_ (.A1(_1313_),
    .A2(_1317_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4798_ (.A1(_1315_),
    .A2(_1176_),
    .B(_1311_),
    .C(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4799_ (.A1(_1315_),
    .A2(_1176_),
    .A3(_1311_),
    .B(_1468_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4800_ (.A1(_1464_),
    .A2(_1466_),
    .A3(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4801_ (.A1(_1459_),
    .A2(_1463_),
    .A3(_1470_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4802_ (.A1(_1454_),
    .A2(_1457_),
    .A3(_1471_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4803_ (.A1(_1444_),
    .A2(_1452_),
    .A3(_1472_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4804_ (.A1(_1406_),
    .A2(_1432_),
    .A3(_1473_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4805_ (.A1(_1328_),
    .A2(_1386_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4806_ (.A1(_1328_),
    .A2(_1386_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4807_ (.A1(_1325_),
    .A2(_1475_),
    .B(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4808_ (.A1(_0625_),
    .A2(_1367_),
    .A3(_1368_),
    .A4(_1381_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4809_ (.A1(_1372_),
    .A2(_1380_),
    .B(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4810_ (.A1(_1365_),
    .A2(_1382_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4811_ (.A1(_1363_),
    .A2(_1383_),
    .B(_1480_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4812_ (.A1(_1477_),
    .A2(_1479_),
    .A3(_1481_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4813_ (.A1(_1399_),
    .A2(_1474_),
    .A3(_1482_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4814_ (.A1(_1396_),
    .A2(_1483_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4815_ (.A1(_1395_),
    .A2(_1392_),
    .A3(_1484_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4816_ (.A1(_1395_),
    .A2(_1392_),
    .B(_1484_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4817_ (.A1(_0803_),
    .A2(_0678_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4818_ (.A1(_0679_),
    .A2(_0680_),
    .A3(\mod.Arithmetic.I_out[79] ),
    .A4(_0681_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4819_ (.A1(_1268_),
    .A2(_1485_),
    .A3(_1486_),
    .B1(_1487_),
    .B2(_1488_),
    .ZN(\mod.P3.Res[7] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4820_ (.I(\mod.Data_Mem.F_M.src[8] ),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4821_ (.I(_1489_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4822_ (.I(_1490_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4823_ (.I(\mod.Data_Mem.F_M.src[1] ),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4824_ (.I(_1492_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4825_ (.I(_1493_),
    .Z(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4826_ (.I(\mod.Data_Mem.F_M.src[2] ),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4827_ (.I(\mod.Data_Mem.F_M.src[4] ),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4828_ (.A1(_1495_),
    .A2(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4829_ (.A1(_1494_),
    .A2(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4830_ (.I(_1498_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4831_ (.I(_1496_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4832_ (.I(\mod.Data_Mem.F_M.src[2] ),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4833_ (.I(_1501_),
    .Z(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4834_ (.I(\mod.Data_Mem.F_M.src[0] ),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4835_ (.I(\mod.Data_Mem.F_M.src[1] ),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4836_ (.A1(_1503_),
    .A2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4837_ (.A1(_1502_),
    .A2(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4838_ (.A1(_1500_),
    .A2(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4839_ (.I(_1507_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4840_ (.I(_1508_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4841_ (.I(_1503_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4842_ (.I(_1510_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4843_ (.I(_1511_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4844_ (.I0(\mod.Data_Mem.F_M.MRAM[21][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][0] ),
    .S(_1512_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4845_ (.I(_1510_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4846_ (.I(_1514_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4847_ (.I0(\mod.Data_Mem.F_M.MRAM[19][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][0] ),
    .S(_1515_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4848_ (.I(_1503_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4849_ (.I(_1517_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4850_ (.I(_1518_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4851_ (.I0(\mod.Data_Mem.F_M.MRAM[17][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][0] ),
    .S(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4852_ (.I(\mod.Data_Mem.F_M.src[0] ),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4853_ (.I(_1521_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4854_ (.A1(_1522_),
    .A2(_1492_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4855_ (.A1(_1505_),
    .A2(_1523_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4856_ (.I(_1524_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4857_ (.I(_1525_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4858_ (.A1(_1521_),
    .A2(_1492_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4859_ (.A1(_1502_),
    .A2(_1527_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4860_ (.I(_1528_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4861_ (.I(_1529_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4862_ (.I0(\mod.Data_Mem.F_M.MRAM[22][0] ),
    .I1(_1513_),
    .I2(_1516_),
    .I3(_1520_),
    .S0(_1526_),
    .S1(_1530_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4863_ (.I(_1497_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4864_ (.I(\mod.Data_Mem.F_M.src[4] ),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4865_ (.I(_1533_),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4866_ (.I(_1534_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4867_ (.I(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4868_ (.I(_1527_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4869_ (.I(_1537_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4870_ (.I(_1538_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4871_ (.I(_1529_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4872_ (.I(\mod.Data_Mem.F_M.src[0] ),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4873_ (.I(_1541_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4874_ (.I(_1542_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4875_ (.I0(\mod.Data_Mem.F_M.MRAM[5][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][0] ),
    .S(_1543_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4876_ (.A1(_1503_),
    .A2(_1504_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4877_ (.I(_1545_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4878_ (.I(_1546_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4879_ (.I0(\mod.Data_Mem.F_M.MRAM[6][0] ),
    .I1(_1544_),
    .S(_1547_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4880_ (.A1(\mod.Data_Mem.F_M.MRAM[3][0] ),
    .A2(_1539_),
    .B1(_1540_),
    .B2(_1548_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4881_ (.A1(_1536_),
    .A2(_1549_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4882_ (.A1(_1509_),
    .A2(_1531_),
    .B(_1532_),
    .C(_1550_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4883_ (.I(\mod.Data_Mem.F_M.src[2] ),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4884_ (.I(_1552_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4885_ (.I(_1505_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4886_ (.A1(_1553_),
    .A2(_1554_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4887_ (.I(_1555_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4888_ (.I(_1556_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4889_ (.A1(_1552_),
    .A2(_1537_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4890_ (.A1(_1534_),
    .A2(_1558_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4891_ (.I(_1559_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4892_ (.I(_1560_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4893_ (.A1(\mod.Data_Mem.F_M.MRAM[15][0] ),
    .A2(_1536_),
    .B1(\mod.Data_Mem.F_M.MRAM[31][0] ),
    .B2(_1561_),
    .C(_1556_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4894_ (.A1(_1551_),
    .A2(_1557_),
    .B(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4895_ (.A1(_1495_),
    .A2(_1505_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4896_ (.I(_1564_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4897_ (.I(_1565_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4898_ (.I(_1524_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4899_ (.I(_1567_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4900_ (.I(_1568_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4901_ (.I(_1543_),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4902_ (.I0(\mod.Data_Mem.F_M.MRAM[773][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][0] ),
    .S(_1570_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4903_ (.A1(_1569_),
    .A2(_1571_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(_1527_),
    .A2(_1545_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4905_ (.I(_1573_),
    .Z(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4906_ (.I(_1574_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4907_ (.I(_1575_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4908_ (.I(_1576_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4909_ (.A1(\mod.Data_Mem.F_M.MRAM[774][0] ),
    .A2(_1577_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4910_ (.A1(_1566_),
    .A2(_1572_),
    .A3(_1578_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4911_ (.I(_1573_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4912_ (.I(_1580_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4913_ (.I(_1581_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4914_ (.I(_1541_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4915_ (.I(_1583_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4916_ (.I(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4917_ (.I0(\mod.Data_Mem.F_M.MRAM[771][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][0] ),
    .S(_1585_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4918_ (.A1(_1582_),
    .A2(_1586_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4919_ (.I(_1567_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4920_ (.I(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4921_ (.I0(\mod.Data_Mem.F_M.MRAM[769][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[768][0] ),
    .S(_1585_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4922_ (.I(_1564_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4923_ (.A1(_1589_),
    .A2(_1590_),
    .B(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4924_ (.A1(_1587_),
    .A2(_1592_),
    .B(_1561_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4925_ (.I(_1492_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4926_ (.A1(_1594_),
    .A2(_1552_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4927_ (.A1(_1518_),
    .A2(_1595_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4928_ (.I(_1596_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4929_ (.I(_1597_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4930_ (.I(_1523_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4931_ (.I(_1599_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4932_ (.I(_1524_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4933_ (.I(_1601_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4934_ (.I(_1517_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4935_ (.I(_1603_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4936_ (.I0(\mod.Data_Mem.F_M.MRAM[789][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][0] ),
    .S(_1604_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4937_ (.A1(\mod.Data_Mem.F_M.MRAM[790][0] ),
    .A2(_1600_),
    .B1(_1602_),
    .B2(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4938_ (.I(_1574_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4939_ (.I(_1607_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4940_ (.I(_1541_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4941_ (.I(_1609_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4942_ (.I(_1610_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4943_ (.I0(\mod.Data_Mem.F_M.MRAM[787][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[786][0] ),
    .S(_1611_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4944_ (.A1(_1608_),
    .A2(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4945_ (.I(_1601_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4946_ (.I(_1603_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4947_ (.I0(\mod.Data_Mem.F_M.MRAM[785][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][0] ),
    .S(_1615_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4948_ (.I(_1564_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4949_ (.A1(_1614_),
    .A2(_1616_),
    .B(_1617_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4950_ (.I(_1507_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4951_ (.A1(_1566_),
    .A2(_1606_),
    .B1(_1613_),
    .B2(_1618_),
    .C(_1619_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4952_ (.A1(_1579_),
    .A2(_1593_),
    .B(_1598_),
    .C(_1620_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4953_ (.I(_1500_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4954_ (.I(_1622_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4955_ (.I(_1508_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4956_ (.A1(_1623_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][0] ),
    .B1(_1624_),
    .B2(\mod.Data_Mem.F_M.MRAM[783][0] ),
    .C(_1556_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4957_ (.A1(_1621_),
    .A2(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4958_ (.A1(_1502_),
    .A2(_1533_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4959_ (.I(_1627_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4960_ (.A1(_1539_),
    .A2(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4961_ (.A1(_1490_),
    .A2(_1629_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4962_ (.A1(_1491_),
    .A2(_1499_),
    .A3(_1563_),
    .B1(_1626_),
    .B2(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4963_ (.I(_1631_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4964_ (.I(_1629_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4965_ (.I(_1622_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4966_ (.I(\mod.Data_Mem.F_M.MRAM[31][1] ),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4967_ (.I(_1619_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4968_ (.A1(_1633_),
    .A2(_1634_),
    .B1(_1635_),
    .B2(\mod.Data_Mem.F_M.MRAM[15][1] ),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4969_ (.I(_1567_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4970_ (.I(_1637_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4971_ (.I(_1603_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4972_ (.I0(\mod.Data_Mem.F_M.MRAM[5][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][1] ),
    .S(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4973_ (.A1(_1638_),
    .A2(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4974_ (.I(_1599_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4975_ (.I(_1642_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4976_ (.I(_1528_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4977_ (.I(_1644_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4978_ (.A1(\mod.Data_Mem.F_M.MRAM[6][1] ),
    .A2(_1643_),
    .B(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4979_ (.I(_1574_),
    .Z(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4980_ (.I(_1647_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4981_ (.I(_1510_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4982_ (.I0(\mod.Data_Mem.F_M.MRAM[3][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][1] ),
    .S(_1649_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4983_ (.I(_1542_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4984_ (.I0(\mod.Data_Mem.F_M.MRAM[1][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][1] ),
    .S(_1651_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4985_ (.A1(_1588_),
    .A2(_1652_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4986_ (.A1(_1648_),
    .A2(_1650_),
    .B(_1653_),
    .C(_1617_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4987_ (.I(_1559_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4988_ (.A1(_1641_),
    .A2(_1646_),
    .B(_1654_),
    .C(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4989_ (.I(_1588_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4990_ (.I(_1603_),
    .Z(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4991_ (.I0(\mod.Data_Mem.F_M.MRAM[17][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][1] ),
    .S(_1658_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4992_ (.A1(_1657_),
    .A2(_1659_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4993_ (.I(_1580_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4994_ (.I(_1661_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4995_ (.I0(\mod.Data_Mem.F_M.MRAM[19][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][1] ),
    .S(_1519_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4996_ (.I(_1564_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4997_ (.A1(_1662_),
    .A2(_1663_),
    .B(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4998_ (.I(_1529_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4999_ (.A1(\mod.Data_Mem.F_M.MRAM[22][1] ),
    .A2(_1643_),
    .B(_1666_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5000_ (.I0(\mod.Data_Mem.F_M.MRAM[21][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][1] ),
    .S(_1639_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5001_ (.A1(_1589_),
    .A2(_1668_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5002_ (.A1(_1660_),
    .A2(_1665_),
    .B1(_1667_),
    .B2(_1669_),
    .C(_1619_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5003_ (.I(_1555_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5004_ (.A1(_1656_),
    .A2(_1670_),
    .B(_1671_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5005_ (.I(\mod.Data_Mem.F_M.src[8] ),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5006_ (.I(_1673_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5007_ (.I(_1674_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5008_ (.I(_1675_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5009_ (.A1(_1557_),
    .A2(_1636_),
    .B(_1672_),
    .C(_1676_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5010_ (.I(_1596_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5011_ (.I(_1678_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5012_ (.I(_1597_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5013_ (.I(_1584_),
    .Z(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5014_ (.I(_1518_),
    .Z(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5015_ (.I(\mod.Data_Mem.F_M.MRAM[784][1] ),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5016_ (.A1(_1682_),
    .A2(_1683_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5017_ (.A1(_1681_),
    .A2(\mod.Data_Mem.F_M.MRAM[785][1] ),
    .B(_1684_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5018_ (.I(\mod.Data_Mem.F_M.MRAM[786][1] ),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5019_ (.A1(_1515_),
    .A2(_1686_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5020_ (.A1(_1681_),
    .A2(\mod.Data_Mem.F_M.MRAM[787][1] ),
    .B(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5021_ (.I(\mod.Data_Mem.F_M.MRAM[788][1] ),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5022_ (.A1(_1570_),
    .A2(_1689_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5023_ (.A1(_1681_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][1] ),
    .B(_1690_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5024_ (.I(_1522_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5025_ (.I(_1692_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5026_ (.I(_1541_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5027_ (.I(_1694_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5028_ (.A1(_1695_),
    .A2(\mod.Data_Mem.F_M.MRAM[790][1] ),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5029_ (.A1(_1693_),
    .A2(\mod.Data_Mem.F_M.MRAM[791][1] ),
    .B(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5030_ (.I(_1575_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5031_ (.I0(_1685_),
    .I1(_1688_),
    .I2(_1691_),
    .I3(_1697_),
    .S0(_1698_),
    .S1(_1565_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5032_ (.A1(_1680_),
    .A2(_1699_),
    .B(_1561_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5033_ (.A1(\mod.Data_Mem.F_M.MRAM[799][1] ),
    .A2(_1679_),
    .B(_1700_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5034_ (.I(_1678_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5035_ (.I(_1565_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5036_ (.I(_1609_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5037_ (.I0(\mod.Data_Mem.F_M.MRAM[773][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][1] ),
    .S(_1704_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5038_ (.I(_1542_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5039_ (.I0(\mod.Data_Mem.F_M.MRAM[775][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][1] ),
    .S(_1706_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5040_ (.I(_1574_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5041_ (.I0(_1705_),
    .I1(_1707_),
    .S(_1708_),
    .Z(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5042_ (.I(_1517_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5043_ (.I(_1710_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5044_ (.I(_1542_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5045_ (.I(\mod.Data_Mem.F_M.MRAM[770][1] ),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5046_ (.A1(_1712_),
    .A2(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5047_ (.A1(_1711_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][1] ),
    .B(_1714_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5048_ (.A1(_1648_),
    .A2(_1715_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5049_ (.I(_1704_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5050_ (.I(_1610_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5051_ (.I(\mod.Data_Mem.F_M.MRAM[768][1] ),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5052_ (.A1(_1718_),
    .A2(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5053_ (.A1(_1717_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][1] ),
    .B(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5054_ (.A1(_1602_),
    .A2(_1721_),
    .B(_1617_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5055_ (.A1(_1703_),
    .A2(_1709_),
    .B1(_1716_),
    .B2(_1722_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5056_ (.I(_1508_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5057_ (.A1(_1680_),
    .A2(_1723_),
    .B(_1724_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5058_ (.A1(\mod.Data_Mem.F_M.MRAM[783][1] ),
    .A2(_1702_),
    .B(_1725_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5059_ (.I(_1673_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5060_ (.I(_1727_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5061_ (.A1(_1701_),
    .A2(_1726_),
    .B(_1728_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5062_ (.A1(_1632_),
    .A2(_1677_),
    .A3(_1729_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5063_ (.I(_1730_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5064_ (.I(_1538_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5065_ (.I(_1567_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5066_ (.I(_1732_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5067_ (.I0(\mod.Data_Mem.F_M.MRAM[5][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][2] ),
    .S(_1639_),
    .Z(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5068_ (.A1(_1733_),
    .A2(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5069_ (.A1(\mod.Data_Mem.F_M.MRAM[6][2] ),
    .A2(_1600_),
    .B(_1644_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5070_ (.I(_1732_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5071_ (.I0(\mod.Data_Mem.F_M.MRAM[1][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][2] ),
    .S(_1519_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5072_ (.A1(_1737_),
    .A2(_1738_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5073_ (.I(_1575_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5074_ (.I0(\mod.Data_Mem.F_M.MRAM[3][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][2] ),
    .S(_1519_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5075_ (.A1(_1740_),
    .A2(_1741_),
    .B(_1617_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5076_ (.A1(_1735_),
    .A2(_1736_),
    .B1(_1739_),
    .B2(_1742_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5077_ (.I0(\mod.Data_Mem.F_M.MRAM[17][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][2] ),
    .S(_1658_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5078_ (.A1(_1602_),
    .A2(_1744_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5079_ (.I(_1607_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5080_ (.I(_1517_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5081_ (.I0(\mod.Data_Mem.F_M.MRAM[19][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][2] ),
    .S(_1747_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5082_ (.A1(_1746_),
    .A2(_1748_),
    .B(_1565_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5083_ (.I(_1599_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5084_ (.A1(\mod.Data_Mem.F_M.MRAM[22][2] ),
    .A2(_1750_),
    .B(_1644_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5085_ (.I(_1601_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5086_ (.I0(\mod.Data_Mem.F_M.MRAM[21][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][2] ),
    .S(_1695_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5087_ (.A1(_1752_),
    .A2(_1753_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5088_ (.A1(_1745_),
    .A2(_1749_),
    .B1(_1751_),
    .B2(_1754_),
    .C(_1619_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5089_ (.A1(_1509_),
    .A2(_1743_),
    .B(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5090_ (.I(_1500_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5091_ (.I(_1757_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5092_ (.A1(_1758_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][2] ),
    .B1(_1724_),
    .B2(\mod.Data_Mem.F_M.MRAM[15][2] ),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5093_ (.I0(_1756_),
    .I1(_1759_),
    .S(_1598_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5094_ (.I(_1674_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5095_ (.I(_1761_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5096_ (.I(_1710_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5097_ (.I0(\mod.Data_Mem.F_M.MRAM[775][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][2] ),
    .S(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5098_ (.I0(\mod.Data_Mem.F_M.MRAM[773][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][2] ),
    .S(_1763_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5099_ (.I0(_1764_),
    .I1(_1765_),
    .S(_1568_),
    .Z(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5100_ (.I(_1704_),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5101_ (.I(_1583_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5102_ (.I(_1768_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5103_ (.I(\mod.Data_Mem.F_M.MRAM[770][2] ),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5104_ (.A1(_1769_),
    .A2(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5105_ (.A1(_1767_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][2] ),
    .B(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5106_ (.A1(_1662_),
    .A2(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5107_ (.I(_1706_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5108_ (.I(\mod.Data_Mem.F_M.MRAM[768][2] ),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5109_ (.A1(_1769_),
    .A2(_1775_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5110_ (.A1(_1774_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][2] ),
    .B(_1776_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5111_ (.A1(_1733_),
    .A2(_1777_),
    .B(_1664_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5112_ (.A1(_1566_),
    .A2(_1766_),
    .B1(_1773_),
    .B2(_1778_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5113_ (.I(_1597_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5114_ (.A1(\mod.Data_Mem.F_M.MRAM[783][2] ),
    .A2(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5115_ (.A1(_1598_),
    .A2(_1779_),
    .B(_1781_),
    .C(_1509_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5116_ (.I(_1692_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5117_ (.A1(_1658_),
    .A2(\mod.Data_Mem.F_M.MRAM[790][2] ),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5118_ (.A1(_1783_),
    .A2(\mod.Data_Mem.F_M.MRAM[791][2] ),
    .B(_1784_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5119_ (.I(_1649_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5120_ (.I(_1609_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5121_ (.I(\mod.Data_Mem.F_M.MRAM[788][2] ),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5122_ (.A1(_1787_),
    .A2(_1788_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5123_ (.A1(_1786_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][2] ),
    .B(_1789_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5124_ (.I(_1706_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5125_ (.I(_1518_),
    .Z(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5126_ (.I(\mod.Data_Mem.F_M.MRAM[786][2] ),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5127_ (.A1(_1792_),
    .A2(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5128_ (.A1(_1791_),
    .A2(\mod.Data_Mem.F_M.MRAM[787][2] ),
    .B(_1794_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5129_ (.I(_1763_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5130_ (.I(\mod.Data_Mem.F_M.MRAM[784][2] ),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5131_ (.A1(_1792_),
    .A2(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5132_ (.A1(_1796_),
    .A2(\mod.Data_Mem.F_M.MRAM[785][2] ),
    .B(_1798_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5133_ (.I0(_1785_),
    .I1(_1790_),
    .I2(_1795_),
    .I3(_1799_),
    .S0(_1526_),
    .S1(_1530_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5134_ (.A1(\mod.Data_Mem.F_M.MRAM[799][2] ),
    .A2(_1780_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5135_ (.A1(_1598_),
    .A2(_1800_),
    .B(_1801_),
    .C(_1561_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5136_ (.A1(_1782_),
    .A2(_1802_),
    .B(_1676_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5137_ (.A1(_1731_),
    .A2(_1628_),
    .B1(_1760_),
    .B2(_1762_),
    .C(_1803_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5138_ (.I(_1580_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5139_ (.I(_1804_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5140_ (.A1(_1674_),
    .A2(_1627_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5141_ (.I(_1761_),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5142_ (.I(_1644_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5143_ (.I(_1651_),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5144_ (.I0(\mod.Data_Mem.F_M.MRAM[21][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][3] ),
    .S(_1809_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5145_ (.A1(\mod.Data_Mem.F_M.MRAM[22][3] ),
    .A2(_1600_),
    .B1(_1614_),
    .B2(_1810_),
    .C(_1508_),
    .ZN(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5146_ (.I0(\mod.Data_Mem.F_M.MRAM[5][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][3] ),
    .S(_1611_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5147_ (.I(_1547_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5148_ (.A1(\mod.Data_Mem.F_M.MRAM[6][3] ),
    .A2(_1608_),
    .B1(_1812_),
    .B2(_1813_),
    .C(_1560_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5149_ (.I(_1504_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5150_ (.I(_1815_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5151_ (.I0(\mod.Data_Mem.F_M.MRAM[3][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[1][3] ),
    .I2(\mod.Data_Mem.F_M.MRAM[0][3] ),
    .I3(\mod.Data_Mem.F_M.MRAM[2][3] ),
    .S0(_1816_),
    .S1(_1787_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5152_ (.I0(\mod.Data_Mem.F_M.MRAM[19][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][3] ),
    .S(_1651_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5153_ (.A1(_1581_),
    .A2(_1818_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5154_ (.I0(\mod.Data_Mem.F_M.MRAM[17][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][3] ),
    .S(_1543_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5155_ (.A1(_1637_),
    .A2(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5156_ (.A1(_1560_),
    .A2(_1819_),
    .A3(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5157_ (.A1(_1655_),
    .A2(_1817_),
    .B(_1822_),
    .C(_1645_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5158_ (.A1(_1808_),
    .A2(_1811_),
    .A3(_1814_),
    .B(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5159_ (.A1(_1807_),
    .A2(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5160_ (.I0(\mod.Data_Mem.F_M.MRAM[785][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][3] ),
    .S(_1769_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5161_ (.A1(_1657_),
    .A2(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5162_ (.I0(\mod.Data_Mem.F_M.MRAM[787][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[786][3] ),
    .S(_1615_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5163_ (.A1(_1662_),
    .A2(_1828_),
    .B(_1664_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5164_ (.I(_1661_),
    .Z(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5165_ (.I(_1768_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5166_ (.I0(\mod.Data_Mem.F_M.MRAM[791][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[790][3] ),
    .S(_1831_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5167_ (.I(_1529_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5168_ (.A1(_1830_),
    .A2(_1832_),
    .B(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5169_ (.I(_1511_),
    .Z(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5170_ (.I0(\mod.Data_Mem.F_M.MRAM[789][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][3] ),
    .S(_1835_),
    .Z(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5171_ (.A1(_1589_),
    .A2(_1836_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5172_ (.A1(_1827_),
    .A2(_1829_),
    .B1(_1834_),
    .B2(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5173_ (.I(_1647_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5174_ (.I(_1692_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5175_ (.A1(_1704_),
    .A2(\mod.Data_Mem.F_M.MRAM[774][3] ),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5176_ (.A1(_1840_),
    .A2(\mod.Data_Mem.F_M.MRAM[775][3] ),
    .B(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5177_ (.A1(_1839_),
    .A2(_1842_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5178_ (.I(_1525_),
    .Z(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5179_ (.I(_1514_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5180_ (.I(\mod.Data_Mem.F_M.MRAM[772][3] ),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5181_ (.A1(_1604_),
    .A2(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5182_ (.A1(_1845_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][3] ),
    .B(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5183_ (.A1(_1844_),
    .A2(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5184_ (.A1(_1591_),
    .A2(_1843_),
    .A3(_1849_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5185_ (.I(\mod.Data_Mem.F_M.MRAM[770][3] ),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5186_ (.A1(_1604_),
    .A2(_1851_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5187_ (.A1(_1845_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][3] ),
    .B(_1852_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5188_ (.A1(_1839_),
    .A2(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5189_ (.I(\mod.Data_Mem.F_M.MRAM[768][3] ),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5190_ (.A1(_1649_),
    .A2(_1855_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5191_ (.A1(_1845_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][3] ),
    .B(_1856_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5192_ (.A1(_1844_),
    .A2(_1857_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5193_ (.A1(_1808_),
    .A2(_1854_),
    .A3(_1858_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5194_ (.A1(_1724_),
    .A2(_1850_),
    .A3(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5195_ (.A1(_1624_),
    .A2(_1838_),
    .B(_1860_),
    .C(_1490_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5196_ (.A1(_1557_),
    .A2(_1825_),
    .A3(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5197_ (.I(_1655_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5198_ (.A1(\mod.Data_Mem.F_M.MRAM[783][3] ),
    .A2(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5199_ (.I(_1489_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5200_ (.A1(\mod.Data_Mem.F_M.MRAM[799][3] ),
    .A2(_1635_),
    .B(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5201_ (.A1(_1758_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][3] ),
    .B1(\mod.Data_Mem.F_M.MRAM[31][3] ),
    .B2(_1724_),
    .C(_1675_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5202_ (.A1(_1864_),
    .A2(_1866_),
    .B(_1867_),
    .C(_1702_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5203_ (.A1(_1632_),
    .A2(_1862_),
    .A3(_1868_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5204_ (.A1(_1805_),
    .A2(_1806_),
    .B(_1869_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5205_ (.I(\mod.Data_Mem.F_M.MRAM[15][4] ),
    .Z(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5206_ (.A1(_1870_),
    .A2(_1679_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5207_ (.I(_1555_),
    .Z(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5208_ (.I(_1583_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5209_ (.I(_1873_),
    .Z(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5210_ (.I0(\mod.Data_Mem.F_M.MRAM[5][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][4] ),
    .S(_1874_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5211_ (.I(_1873_),
    .Z(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5212_ (.I0(\mod.Data_Mem.F_M.MRAM[7][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][4] ),
    .S(_1876_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5213_ (.I(_1584_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5214_ (.I0(\mod.Data_Mem.F_M.MRAM[1][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][4] ),
    .S(_1878_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5215_ (.I(_1873_),
    .Z(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5216_ (.I0(\mod.Data_Mem.F_M.MRAM[3][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][4] ),
    .S(_1880_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5217_ (.I(_1647_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5218_ (.I0(_1875_),
    .I1(_1877_),
    .I2(_1879_),
    .I3(_1881_),
    .S0(_1882_),
    .S1(_1666_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5219_ (.I(_1560_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5220_ (.A1(_1872_),
    .A2(_1883_),
    .B(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5221_ (.I(_1678_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5222_ (.A1(\mod.Data_Mem.F_M.MRAM[31][4] ),
    .A2(_1886_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5223_ (.I(_1555_),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5224_ (.I(_1609_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5225_ (.I(_1889_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5226_ (.I0(\mod.Data_Mem.F_M.MRAM[23][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][4] ),
    .S(_1890_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5227_ (.I(_1610_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5228_ (.I0(\mod.Data_Mem.F_M.MRAM[21][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][4] ),
    .S(_1892_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5229_ (.I0(\mod.Data_Mem.F_M.MRAM[19][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][4] ),
    .S(_1718_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5230_ (.I0(\mod.Data_Mem.F_M.MRAM[17][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][4] ),
    .S(_1718_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5231_ (.I(_1601_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5232_ (.I0(_1891_),
    .I1(_1893_),
    .I2(_1894_),
    .I3(_1895_),
    .S0(_1896_),
    .S1(_1666_),
    .Z(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5233_ (.A1(_1888_),
    .A2(_1897_),
    .B(_1635_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5234_ (.I(_1674_),
    .Z(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5235_ (.A1(_1899_),
    .A2(_1629_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5236_ (.A1(_1871_),
    .A2(_1885_),
    .B1(_1887_),
    .B2(_1898_),
    .C(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5237_ (.I(\mod.Data_Mem.F_M.MRAM[783][4] ),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5238_ (.A1(_1902_),
    .A2(_1702_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5239_ (.I(_1514_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5240_ (.I0(\mod.Data_Mem.F_M.MRAM[773][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][4] ),
    .S(_1904_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5241_ (.I(_1768_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5242_ (.I0(\mod.Data_Mem.F_M.MRAM[775][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][4] ),
    .S(_1906_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5243_ (.I(_1514_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5244_ (.I0(\mod.Data_Mem.F_M.MRAM[769][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[768][4] ),
    .S(_1908_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5245_ (.I0(\mod.Data_Mem.F_M.MRAM[771][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][4] ),
    .S(_1831_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5246_ (.I(_1647_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5247_ (.I0(_1905_),
    .I1(_1907_),
    .I2(_1909_),
    .I3(_1910_),
    .S0(_1911_),
    .S1(_1645_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5248_ (.A1(_1557_),
    .A2(_1912_),
    .B(_1863_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5249_ (.I(_1678_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5250_ (.I(_1543_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5251_ (.I(_1504_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5252_ (.I(_1916_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5253_ (.I0(\mod.Data_Mem.F_M.MRAM[791][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][4] ),
    .I2(\mod.Data_Mem.F_M.MRAM[789][4] ),
    .I3(\mod.Data_Mem.F_M.MRAM[790][4] ),
    .S0(_1915_),
    .S1(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5254_ (.A1(_1703_),
    .A2(_1918_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5255_ (.I(_1732_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5256_ (.I(_1694_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5257_ (.I(\mod.Data_Mem.F_M.MRAM[787][4] ),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5258_ (.I(_1694_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5259_ (.A1(_1923_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][4] ),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5260_ (.A1(_1921_),
    .A2(_1922_),
    .B(_1924_),
    .ZN(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5261_ (.I0(\mod.Data_Mem.F_M.MRAM[785][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][4] ),
    .S(_1610_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5262_ (.A1(_1576_),
    .A2(_1926_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5263_ (.A1(_1920_),
    .A2(_1925_),
    .B(_1927_),
    .C(_1833_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5264_ (.A1(_1919_),
    .A2(_1928_),
    .B(_1680_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5265_ (.A1(\mod.Data_Mem.F_M.MRAM[799][4] ),
    .A2(_1914_),
    .B(_1929_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5266_ (.I(_1655_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5267_ (.A1(_1903_),
    .A2(_1913_),
    .B1(_1930_),
    .B2(_1931_),
    .C(_1630_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5268_ (.A1(_1901_),
    .A2(_1932_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5269_ (.I(_1933_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5270_ (.I(_1597_),
    .Z(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5271_ (.A1(\mod.Data_Mem.F_M.MRAM[799][5] ),
    .A2(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5272_ (.I(_1698_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5273_ (.I(_1889_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5274_ (.I(\mod.Data_Mem.F_M.MRAM[788][5] ),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5275_ (.A1(_1921_),
    .A2(_1938_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5276_ (.A1(_1937_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][5] ),
    .B(_1939_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5277_ (.I0(\mod.Data_Mem.F_M.MRAM[791][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[790][5] ),
    .S(_1512_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5278_ (.A1(_1830_),
    .A2(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5279_ (.A1(_1936_),
    .A2(_1940_),
    .B(_1942_),
    .C(_1566_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5280_ (.I(_1583_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5281_ (.I0(\mod.Data_Mem.F_M.MRAM[787][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[786][5] ),
    .S(_1944_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5282_ (.A1(_1582_),
    .A2(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5283_ (.I0(\mod.Data_Mem.F_M.MRAM[785][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][5] ),
    .S(_1874_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5284_ (.A1(_1569_),
    .A2(_1947_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5285_ (.A1(_1808_),
    .A2(_1946_),
    .A3(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5286_ (.A1(_1671_),
    .A2(_1943_),
    .A3(_1949_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5287_ (.A1(_1931_),
    .A2(_1935_),
    .A3(_1950_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5288_ (.I0(\mod.Data_Mem.F_M.MRAM[773][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][5] ),
    .S(_1876_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5289_ (.I0(\mod.Data_Mem.F_M.MRAM[775][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][5] ),
    .S(_1585_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5290_ (.I(_1710_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5291_ (.I(\mod.Data_Mem.F_M.MRAM[769][5] ),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5292_ (.I(_1651_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5293_ (.A1(_1956_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][5] ),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5294_ (.A1(_1954_),
    .A2(_1955_),
    .B(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5295_ (.I0(\mod.Data_Mem.F_M.MRAM[771][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][5] ),
    .S(_1874_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5296_ (.I0(_1952_),
    .I1(_1953_),
    .I2(_1958_),
    .I3(_1959_),
    .S0(_1882_),
    .S1(_1645_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5297_ (.A1(_1888_),
    .A2(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5298_ (.A1(\mod.Data_Mem.F_M.MRAM[783][5] ),
    .A2(_1934_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5299_ (.A1(_1635_),
    .A2(_1961_),
    .A3(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5300_ (.A1(_1632_),
    .A2(_1951_),
    .A3(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5301_ (.A1(\mod.Data_Mem.F_M.MRAM[15][5] ),
    .A2(_1934_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5302_ (.I0(\mod.Data_Mem.F_M.MRAM[5][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][5] ),
    .S(_1570_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5303_ (.I0(\mod.Data_Mem.F_M.MRAM[7][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][5] ),
    .S(_1682_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5304_ (.I(\mod.Data_Mem.F_M.MRAM[1][5] ),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5305_ (.A1(_1906_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][5] ),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5306_ (.A1(_1711_),
    .A2(_1968_),
    .B(_1969_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5307_ (.I(_1511_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5308_ (.I0(\mod.Data_Mem.F_M.MRAM[3][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][5] ),
    .S(_1971_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5309_ (.I0(_1966_),
    .I1(_1967_),
    .I2(_1970_),
    .I3(_1972_),
    .S0(_1698_),
    .S1(_1530_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5310_ (.A1(_1671_),
    .A2(_1973_),
    .B(_1884_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5311_ (.A1(\mod.Data_Mem.F_M.MRAM[31][5] ),
    .A2(_1934_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5312_ (.I0(\mod.Data_Mem.F_M.MRAM[23][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][5] ),
    .S(_1971_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5313_ (.I0(\mod.Data_Mem.F_M.MRAM[21][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][5] ),
    .S(_1570_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5314_ (.I0(\mod.Data_Mem.F_M.MRAM[19][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][5] ),
    .S(_1604_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5315_ (.I0(\mod.Data_Mem.F_M.MRAM[17][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][5] ),
    .S(_1971_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5316_ (.I0(_1976_),
    .I1(_1977_),
    .I2(_1978_),
    .I3(_1979_),
    .S0(_1526_),
    .S1(_1530_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5317_ (.A1(_1556_),
    .A2(_1980_),
    .B(_1509_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5318_ (.A1(_1965_),
    .A2(_1974_),
    .B1(_1975_),
    .B2(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5319_ (.A1(_1491_),
    .A2(_1982_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5320_ (.A1(_1900_),
    .A2(_1964_),
    .B(_1983_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5321_ (.A1(\mod.Data_Mem.F_M.MRAM[15][6] ),
    .A2(_1679_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5322_ (.I0(\mod.Data_Mem.F_M.MRAM[5][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][6] ),
    .S(_1874_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5323_ (.I0(\mod.Data_Mem.F_M.MRAM[7][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][6] ),
    .S(_1876_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5324_ (.I0(\mod.Data_Mem.F_M.MRAM[1][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][6] ),
    .S(_1878_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5325_ (.I0(\mod.Data_Mem.F_M.MRAM[3][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][6] ),
    .S(_1890_),
    .Z(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5326_ (.I0(_1985_),
    .I1(_1986_),
    .I2(_1987_),
    .I3(_1988_),
    .S0(_1882_),
    .S1(_1666_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5327_ (.A1(_1872_),
    .A2(_1989_),
    .B(_1884_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5328_ (.A1(\mod.Data_Mem.F_M.MRAM[31][6] ),
    .A2(_1886_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5329_ (.I0(\mod.Data_Mem.F_M.MRAM[23][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][6] ),
    .S(_1890_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5330_ (.I0(\mod.Data_Mem.F_M.MRAM[21][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][6] ),
    .S(_1892_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5331_ (.I0(\mod.Data_Mem.F_M.MRAM[19][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][6] ),
    .S(_1809_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5332_ (.I0(\mod.Data_Mem.F_M.MRAM[17][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][6] ),
    .S(_1718_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5333_ (.I0(_1992_),
    .I1(_1993_),
    .I2(_1994_),
    .I3(_1995_),
    .S0(_1896_),
    .S1(_1540_),
    .Z(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5334_ (.A1(_1888_),
    .A2(_1996_),
    .B(_1624_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5335_ (.A1(_1984_),
    .A2(_1990_),
    .B1(_1991_),
    .B2(_1997_),
    .C(_1900_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5336_ (.A1(\mod.Data_Mem.F_M.MRAM[783][6] ),
    .A2(_1702_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5337_ (.I0(\mod.Data_Mem.F_M.MRAM[769][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[768][6] ),
    .S(_1904_),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5338_ (.I0(\mod.Data_Mem.F_M.MRAM[771][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][6] ),
    .S(_1906_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5339_ (.I0(\mod.Data_Mem.F_M.MRAM[773][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][6] ),
    .S(_1908_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5340_ (.I0(\mod.Data_Mem.F_M.MRAM[775][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][6] ),
    .S(_1831_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5341_ (.I0(_2000_),
    .I1(_2001_),
    .I2(_2002_),
    .I3(_2003_),
    .S0(_1911_),
    .S1(_1591_),
    .Z(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5342_ (.A1(_1872_),
    .A2(_2004_),
    .B(_1863_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5343_ (.I0(\mod.Data_Mem.F_M.MRAM[791][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][6] ),
    .I2(\mod.Data_Mem.F_M.MRAM[789][6] ),
    .I3(\mod.Data_Mem.F_M.MRAM[790][6] ),
    .S0(_1915_),
    .S1(_1917_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5344_ (.A1(_1703_),
    .A2(_2006_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5345_ (.I(_1732_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5346_ (.I(\mod.Data_Mem.F_M.MRAM[787][6] ),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5347_ (.A1(_1923_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][6] ),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5348_ (.A1(_1921_),
    .A2(_2009_),
    .B(_2010_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5349_ (.I0(\mod.Data_Mem.F_M.MRAM[785][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][6] ),
    .S(_1889_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5350_ (.A1(_1576_),
    .A2(_2012_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5351_ (.A1(_2008_),
    .A2(_2011_),
    .B(_2013_),
    .C(_1833_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5352_ (.A1(_2007_),
    .A2(_2014_),
    .B(_1780_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5353_ (.A1(\mod.Data_Mem.F_M.MRAM[799][6] ),
    .A2(_1914_),
    .B(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5354_ (.A1(_1999_),
    .A2(_2005_),
    .B1(_2016_),
    .B2(_1931_),
    .C(_1630_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5355_ (.A1(_1998_),
    .A2(_2017_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5356_ (.I(_2018_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5357_ (.A1(\mod.Data_Mem.F_M.MRAM[15][7] ),
    .A2(_1886_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5358_ (.I0(\mod.Data_Mem.F_M.MRAM[1][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[0][7] ),
    .S(_1892_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5359_ (.I0(\mod.Data_Mem.F_M.MRAM[3][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][7] ),
    .S(_1876_),
    .Z(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5360_ (.I0(\mod.Data_Mem.F_M.MRAM[5][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[4][7] ),
    .S(_1878_),
    .Z(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5361_ (.I0(\mod.Data_Mem.F_M.MRAM[7][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][7] ),
    .S(_1890_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5362_ (.I0(_2020_),
    .I1(_2021_),
    .I2(_2022_),
    .I3(_2023_),
    .S0(_1698_),
    .S1(_1664_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5363_ (.A1(_1888_),
    .A2(_2024_),
    .B(_1884_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5364_ (.A1(\mod.Data_Mem.F_M.MRAM[31][7] ),
    .A2(_1914_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5365_ (.I0(\mod.Data_Mem.F_M.MRAM[23][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][7] ),
    .S(_1878_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5366_ (.I0(\mod.Data_Mem.F_M.MRAM[21][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[20][7] ),
    .S(_1880_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5367_ (.I0(\mod.Data_Mem.F_M.MRAM[19][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[18][7] ),
    .S(_1809_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5368_ (.I0(\mod.Data_Mem.F_M.MRAM[17][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[16][7] ),
    .S(_1611_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5369_ (.I0(_2027_),
    .I1(_2028_),
    .I2(_2029_),
    .I3(_2030_),
    .S0(_1896_),
    .S1(_1540_),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5370_ (.A1(_1671_),
    .A2(_2031_),
    .B(_1624_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5371_ (.A1(_2019_),
    .A2(_2025_),
    .B1(_2026_),
    .B2(_2032_),
    .C(_1900_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5372_ (.A1(\mod.Data_Mem.F_M.MRAM[783][7] ),
    .A2(_1679_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5373_ (.I0(\mod.Data_Mem.F_M.MRAM[769][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[768][7] ),
    .S(_1904_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5374_ (.I0(\mod.Data_Mem.F_M.MRAM[771][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[770][7] ),
    .S(_1906_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5375_ (.I0(\mod.Data_Mem.F_M.MRAM[773][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[772][7] ),
    .S(_1908_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5376_ (.I0(\mod.Data_Mem.F_M.MRAM[775][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[774][7] ),
    .S(_1831_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5377_ (.I0(_2035_),
    .I1(_2036_),
    .I2(_2037_),
    .I3(_2038_),
    .S0(_1911_),
    .S1(_1591_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5378_ (.A1(_1872_),
    .A2(_2039_),
    .B(_1863_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5379_ (.I0(\mod.Data_Mem.F_M.MRAM[791][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[788][7] ),
    .I2(\mod.Data_Mem.F_M.MRAM[789][7] ),
    .I3(\mod.Data_Mem.F_M.MRAM[790][7] ),
    .S0(_1915_),
    .S1(_1917_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5380_ (.A1(_1703_),
    .A2(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5381_ (.I(\mod.Data_Mem.F_M.MRAM[787][7] ),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5382_ (.A1(_1923_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][7] ),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5383_ (.A1(_1767_),
    .A2(_2043_),
    .B(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5384_ (.I0(\mod.Data_Mem.F_M.MRAM[785][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[784][7] ),
    .S(_1889_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5385_ (.A1(_1576_),
    .A2(_2046_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5386_ (.A1(_2008_),
    .A2(_2045_),
    .B(_2047_),
    .C(_1833_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5387_ (.A1(_2042_),
    .A2(_2048_),
    .B(_1780_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5388_ (.A1(\mod.Data_Mem.F_M.MRAM[799][7] ),
    .A2(_1914_),
    .B(_2049_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5389_ (.A1(_2034_),
    .A2(_2040_),
    .B1(_2050_),
    .B2(_1931_),
    .C(_1630_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5390_ (.A1(_2033_),
    .A2(_2051_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5391_ (.I(_2052_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5392_ (.I(_1522_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5393_ (.I(_2053_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5394_ (.I(_2054_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5395_ (.I(_2055_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5396_ (.I(_2056_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5397_ (.I(_1502_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5398_ (.A1(_2058_),
    .A2(_1534_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5399_ (.A1(_1673_),
    .A2(_2059_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5400_ (.I(_2060_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5401_ (.I(_2061_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5402_ (.I(_2062_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5403_ (.A1(_2057_),
    .A2(_0010_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5404_ (.I(_1594_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5405_ (.I(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5406_ (.I(_2064_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5407_ (.I(_2065_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5408_ (.I(_1727_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5409_ (.I(_2067_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5410_ (.I(_2059_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5411_ (.I(_2069_),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5412_ (.I(_2070_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5413_ (.A1(_2066_),
    .A2(_2068_),
    .A3(_2071_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5414_ (.I(_1673_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5415_ (.I(_2072_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5416_ (.I(_2073_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5417_ (.A1(_2074_),
    .A2(_2071_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5418_ (.I(_1511_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5419_ (.I(_2075_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5420_ (.A1(_2076_),
    .A2(_0010_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5421_ (.I(_2061_),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5422_ (.A1(_1805_),
    .A2(_2077_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5423_ (.I(_2078_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5424_ (.I(\mod.Data_Mem.F_M.src[8] ),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5425_ (.I(_2079_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5426_ (.I(_2080_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5427_ (.I(_1554_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5428_ (.I(_2082_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5429_ (.A1(_2081_),
    .A2(_2083_),
    .A3(_2070_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5430_ (.A1(_2074_),
    .A2(_2071_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5431_ (.A1(_2057_),
    .A2(_0010_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5432_ (.I(_1493_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5433_ (.I(_2084_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5434_ (.A1(_2085_),
    .A2(_2061_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5435_ (.I(_2086_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5436_ (.A1(_2066_),
    .A2(_2068_),
    .A3(_2070_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5437_ (.A1(_2074_),
    .A2(_2071_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5438_ (.I(_1815_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5439_ (.I(_2087_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5440_ (.I(_2088_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5441_ (.I(_1553_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5442_ (.A1(_2090_),
    .A2(_1622_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5443_ (.A1(_1727_),
    .A2(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5444_ (.A1(_2089_),
    .A2(_2092_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5445_ (.I(_1522_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5446_ (.I(_2094_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5447_ (.A1(_1908_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][0] ),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5448_ (.A1(_2095_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][0] ),
    .B(_2096_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5449_ (.I(_1535_),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5450_ (.A1(_1916_),
    .A2(_1495_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5451_ (.I(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5452_ (.I(_2100_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5453_ (.A1(_2098_),
    .A2(_2101_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5454_ (.A1(_2076_),
    .A2(_2102_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5455_ (.I(_1496_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5456_ (.I(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5457_ (.I(_2105_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5458_ (.A1(_2063_),
    .A2(_2058_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5459_ (.I(_2107_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5460_ (.A1(_2106_),
    .A2(_2108_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5461_ (.I0(\mod.Data_Mem.F_M.MRAM[30][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[31][0] ),
    .S(_1712_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5462_ (.I(_1806_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5463_ (.A1(_2111_),
    .A2(_2060_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5464_ (.A1(_2109_),
    .A2(_2110_),
    .B(_2112_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5465_ (.A1(_2093_),
    .A2(_2097_),
    .B1(_2103_),
    .B2(_2113_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5466_ (.I(_1916_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5467_ (.I(_2114_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5468_ (.A1(_2115_),
    .A2(_1627_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5469_ (.I(_2116_),
    .Z(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5470_ (.I(_2086_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5471_ (.A1(_1585_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][1] ),
    .Z(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5472_ (.A1(_2095_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][1] ),
    .B(_2119_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5473_ (.I0(\mod.Data_Mem.F_M.MRAM[798][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[799][1] ),
    .S(_1880_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5474_ (.A1(_2093_),
    .A2(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5475_ (.A1(_2068_),
    .A2(_2117_),
    .B1(_2118_),
    .B2(_2120_),
    .C(_2122_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5476_ (.I0(\mod.Data_Mem.F_M.MRAM[30][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[31][2] ),
    .S(_1682_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5477_ (.I0(\mod.Data_Mem.F_M.MRAM[798][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[799][2] ),
    .S(_1892_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5478_ (.A1(_0025_),
    .A2(_2123_),
    .B1(_2124_),
    .B2(_2093_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5479_ (.A1(_1806_),
    .A2(_2125_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5480_ (.I0(\mod.Data_Mem.F_M.MRAM[30][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[31][3] ),
    .S(_1787_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5481_ (.A1(_2108_),
    .A2(_2126_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5482_ (.I(_2094_),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5483_ (.A1(_1792_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][3] ),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5484_ (.A1(_2128_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][3] ),
    .B(_2129_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5485_ (.A1(_1761_),
    .A2(_2069_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5486_ (.A1(_2066_),
    .A2(_2131_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5487_ (.A1(_2112_),
    .A2(_2127_),
    .B1(_2130_),
    .B2(_2132_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5488_ (.I(_1840_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5489_ (.A1(_1796_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][4] ),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5490_ (.A1(_2133_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][4] ),
    .B(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5491_ (.I(_1692_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5492_ (.A1(_1615_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][4] ),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5493_ (.A1(_2136_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][4] ),
    .B(_2137_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5494_ (.A1(_2118_),
    .A2(_2135_),
    .B1(_2138_),
    .B2(_2132_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5495_ (.A1(_1658_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][5] ),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5496_ (.A1(_1693_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][5] ),
    .B(_2139_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5497_ (.A1(_1835_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][5] ),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5498_ (.I(_2053_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5499_ (.A1(_2142_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][5] ),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5500_ (.A1(_2141_),
    .A2(_2143_),
    .B(_2067_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5501_ (.A1(_2081_),
    .A2(_2140_),
    .B(_2144_),
    .C(_2102_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5502_ (.A1(_1791_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][6] ),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5503_ (.A1(_2133_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][6] ),
    .B(_2145_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5504_ (.A1(_1615_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][6] ),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5505_ (.A1(_1783_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][6] ),
    .B(_2147_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5506_ (.A1(_2118_),
    .A2(_2146_),
    .B1(_2148_),
    .B2(_2132_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5507_ (.A1(_1767_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][7] ),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5508_ (.A1(_2133_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][7] ),
    .B(_2149_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5509_ (.A1(_1809_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][7] ),
    .Z(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5510_ (.A1(_2136_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][7] ),
    .B(_2151_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5511_ (.A1(_2118_),
    .A2(_2150_),
    .B1(_2152_),
    .B2(_2132_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5512_ (.I(_1547_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5513_ (.I(_2153_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5514_ (.A1(_2154_),
    .A2(_2091_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5515_ (.I(_1526_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5516_ (.I(_1682_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5517_ (.I(_2114_),
    .Z(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5518_ (.A1(_2157_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[31][0] ),
    .B2(_2158_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5519_ (.I(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5520_ (.A1(\mod.Data_Mem.F_M.MRAM[29][0] ),
    .A2(_2083_),
    .B1(_2156_),
    .B2(_2160_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5521_ (.I(_2112_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5522_ (.A1(_2076_),
    .A2(_2061_),
    .B1(_2155_),
    .B2(_2161_),
    .C(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5523_ (.I(_2131_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5524_ (.I(_1844_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5525_ (.I(_1815_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5526_ (.I(_2166_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5527_ (.I(_2167_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5528_ (.I(_1711_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5529_ (.A1(_2168_),
    .A2(\mod.Data_Mem.F_M.MRAM[798][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[799][0] ),
    .B2(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5530_ (.A1(_2165_),
    .A2(_2170_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5531_ (.A1(\mod.Data_Mem.F_M.MRAM[797][0] ),
    .A2(_1731_),
    .B(_2171_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5532_ (.A1(_2154_),
    .A2(_2164_),
    .A3(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5533_ (.A1(_2163_),
    .A2(_2173_),
    .Z(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5534_ (.I(_2174_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5535_ (.A1(_2154_),
    .A2(_2131_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5536_ (.I(_2082_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5537_ (.I(_1642_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5538_ (.I(_1575_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5539_ (.I(_1695_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5540_ (.A1(_2179_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][1] ),
    .B2(_1917_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5541_ (.A1(_2178_),
    .A2(_2180_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5542_ (.A1(\mod.Data_Mem.F_M.MRAM[797][1] ),
    .A2(_2176_),
    .B1(_2177_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][1] ),
    .C(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5543_ (.I(_1532_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5544_ (.A1(_2088_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][1] ),
    .B1(_1634_),
    .B2(_1954_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5545_ (.A1(_2008_),
    .A2(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5546_ (.A1(\mod.Data_Mem.F_M.MRAM[29][1] ),
    .A2(_1539_),
    .B1(_1813_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][1] ),
    .C(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5547_ (.A1(_2165_),
    .A2(_2183_),
    .B1(_2155_),
    .B2(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5548_ (.A1(_1762_),
    .A2(_2187_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5549_ (.A1(_2175_),
    .A2(_2182_),
    .B(_2188_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5550_ (.I(_1642_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5551_ (.A1(_1954_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][2] ),
    .B2(_2088_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5552_ (.A1(_1648_),
    .A2(_2190_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5553_ (.A1(\mod.Data_Mem.F_M.MRAM[797][2] ),
    .A2(_2176_),
    .B1(_2189_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][2] ),
    .C(_2191_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5554_ (.I(_1538_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5555_ (.I(_1546_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5556_ (.I(_2194_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5557_ (.I(_2094_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5558_ (.A1(_2064_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[31][2] ),
    .B2(_2196_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5559_ (.A1(_1657_),
    .A2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5560_ (.A1(\mod.Data_Mem.F_M.MRAM[29][2] ),
    .A2(_2193_),
    .B1(_2195_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][2] ),
    .C(_2198_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5561_ (.A1(_2155_),
    .A2(_2199_),
    .B(_1632_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5562_ (.A1(_1762_),
    .A2(_2200_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5563_ (.A1(_2175_),
    .A2(_2192_),
    .B(_2201_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5564_ (.I(_1553_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5565_ (.I(_2202_),
    .Z(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5566_ (.I(_2203_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5567_ (.I(_1600_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5568_ (.I(\mod.Data_Mem.F_M.MRAM[29][3] ),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5569_ (.I(_2054_),
    .Z(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5570_ (.A1(_2207_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][3] ),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5571_ (.I(_2054_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5572_ (.I(_2063_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5573_ (.A1(_2209_),
    .A2(\mod.Data_Mem.F_M.MRAM[30][3] ),
    .B(_2210_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5574_ (.A1(_2206_),
    .A2(_2176_),
    .B1(_2208_),
    .B2(_2211_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5575_ (.A1(_2204_),
    .A2(_2205_),
    .A3(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5576_ (.I(_1554_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5577_ (.A1(_1783_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][3] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][3] ),
    .B2(_2084_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5578_ (.A1(_2214_),
    .A2(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5579_ (.A1(\mod.Data_Mem.F_M.MRAM[797][3] ),
    .A2(_2176_),
    .B1(_2189_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][3] ),
    .C(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5580_ (.I(_2175_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5581_ (.A1(_2112_),
    .A2(_2213_),
    .B1(_2217_),
    .B2(_2218_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5582_ (.I(_1761_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5583_ (.A1(_2219_),
    .A2(_2154_),
    .A3(_2091_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5584_ (.I(_1554_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5585_ (.I(_1599_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5586_ (.I(_1580_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5587_ (.I(_1510_),
    .Z(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5588_ (.I(_1815_),
    .Z(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5589_ (.A1(_2224_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][4] ),
    .B1(\mod.Data_Mem.F_M.MRAM[30][4] ),
    .B2(_2225_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5590_ (.A1(_2223_),
    .A2(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5591_ (.A1(\mod.Data_Mem.F_M.MRAM[29][4] ),
    .A2(_2221_),
    .B1(_2222_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][4] ),
    .C(_2227_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5592_ (.I(_1694_),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5593_ (.A1(_2229_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][4] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][4] ),
    .B2(_1816_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5594_ (.A1(_1708_),
    .A2(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5595_ (.A1(\mod.Data_Mem.F_M.MRAM[797][4] ),
    .A2(_2214_),
    .B1(_1750_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][4] ),
    .C(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5596_ (.A1(_2220_),
    .A2(_2228_),
    .B1(_2232_),
    .B2(_2218_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5597_ (.A1(_2224_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][5] ),
    .B1(\mod.Data_Mem.F_M.MRAM[30][5] ),
    .B2(_2225_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5598_ (.A1(_2223_),
    .A2(_2233_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5599_ (.A1(\mod.Data_Mem.F_M.MRAM[29][5] ),
    .A2(_2221_),
    .B1(_2222_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][5] ),
    .C(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5600_ (.A1(_2229_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][5] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][5] ),
    .B2(_1816_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5601_ (.A1(_1708_),
    .A2(_2236_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5602_ (.A1(\mod.Data_Mem.F_M.MRAM[797][5] ),
    .A2(_2214_),
    .B1(_1750_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][5] ),
    .C(_2237_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5603_ (.A1(_2220_),
    .A2(_2235_),
    .B1(_2238_),
    .B2(_2218_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5604_ (.A1(_1747_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][6] ),
    .B1(\mod.Data_Mem.F_M.MRAM[30][6] ),
    .B2(_2166_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5605_ (.A1(_2223_),
    .A2(_2239_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5606_ (.A1(\mod.Data_Mem.F_M.MRAM[29][6] ),
    .A2(_2082_),
    .B1(_2222_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][6] ),
    .C(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5607_ (.A1(_2229_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][6] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][6] ),
    .B2(_1816_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5608_ (.A1(_1708_),
    .A2(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5609_ (.A1(\mod.Data_Mem.F_M.MRAM[797][6] ),
    .A2(_2221_),
    .B1(_1750_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][6] ),
    .C(_2243_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5610_ (.A1(_2220_),
    .A2(_2241_),
    .B1(_2244_),
    .B2(_2218_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5611_ (.A1(_1747_),
    .A2(\mod.Data_Mem.F_M.MRAM[31][7] ),
    .B1(\mod.Data_Mem.F_M.MRAM[30][7] ),
    .B2(_2166_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5612_ (.A1(_1661_),
    .A2(_2245_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5613_ (.A1(\mod.Data_Mem.F_M.MRAM[29][7] ),
    .A2(_2082_),
    .B1(_1642_),
    .B2(\mod.Data_Mem.F_M.MRAM[28][7] ),
    .C(_2246_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5614_ (.A1(_2229_),
    .A2(\mod.Data_Mem.F_M.MRAM[799][7] ),
    .B1(\mod.Data_Mem.F_M.MRAM[798][7] ),
    .B2(_2225_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5615_ (.A1(_2223_),
    .A2(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5616_ (.A1(\mod.Data_Mem.F_M.MRAM[797][7] ),
    .A2(_2221_),
    .B1(_2222_),
    .B2(\mod.Data_Mem.F_M.MRAM[796][7] ),
    .C(_2249_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5617_ (.A1(_2220_),
    .A2(_2247_),
    .B1(_2250_),
    .B2(_2175_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5618_ (.A1(_2055_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][0] ),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5619_ (.I(_1956_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5620_ (.I(_1493_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5621_ (.I(_2253_),
    .Z(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5622_ (.A1(_2252_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][0] ),
    .B(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5623_ (.A1(_2085_),
    .A2(_2097_),
    .B1(_2251_),
    .B2(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5624_ (.A1(_2092_),
    .A2(_2256_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5625_ (.I(_2069_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5626_ (.I(_2142_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5627_ (.A1(_2259_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][0] ),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5628_ (.I(_1956_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5629_ (.I(_1494_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5630_ (.A1(_2261_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][0] ),
    .B(_2262_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5631_ (.I(_2087_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5632_ (.A1(_2264_),
    .A2(_2110_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5633_ (.A1(_2260_),
    .A2(_2263_),
    .B(_2265_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5634_ (.A1(_2067_),
    .A2(_2258_),
    .A3(_2266_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5635_ (.A1(_2057_),
    .A2(_2111_),
    .B(_2257_),
    .C(_2267_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5636_ (.I(_2053_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5637_ (.I(_2268_),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5638_ (.A1(_2269_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][1] ),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5639_ (.I(_1706_),
    .Z(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5640_ (.A1(_2271_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][1] ),
    .B(_2262_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5641_ (.I(_1916_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5642_ (.A1(_2273_),
    .A2(_2121_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5643_ (.A1(_2270_),
    .A2(_2272_),
    .B(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5644_ (.A1(_2164_),
    .A2(_2275_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5645_ (.I(_1494_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5646_ (.I(_2094_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5647_ (.A1(_2278_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][1] ),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5648_ (.I(_2063_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5649_ (.A1(_2157_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][1] ),
    .B(_2280_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5650_ (.A1(_2277_),
    .A2(_2120_),
    .B1(_2279_),
    .B2(_2281_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5651_ (.A1(_2062_),
    .A2(_2282_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5652_ (.A1(_2089_),
    .A2(_1806_),
    .B(_2276_),
    .C(_2283_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5653_ (.A1(_2269_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][2] ),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5654_ (.A1(_2271_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][2] ),
    .B(_2262_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5655_ (.A1(_2264_),
    .A2(_2124_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5656_ (.A1(_2284_),
    .A2(_2285_),
    .B(_2286_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(_2164_),
    .A2(_2287_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5658_ (.I(_2054_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5659_ (.A1(_2289_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][2] ),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5660_ (.A1(_2252_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][2] ),
    .B(_2254_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5661_ (.A1(_2273_),
    .A2(_2123_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5662_ (.A1(_2290_),
    .A2(_2291_),
    .B(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5663_ (.A1(_2062_),
    .A2(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5664_ (.A1(_2068_),
    .A2(_2117_),
    .B(_2288_),
    .C(_2294_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5665_ (.A1(_2264_),
    .A2(_2126_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5666_ (.I(_1787_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5667_ (.I(_1611_),
    .Z(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5668_ (.A1(_2297_),
    .A2(_2206_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5669_ (.A1(_2296_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][3] ),
    .B(_2298_),
    .C(_2262_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5670_ (.A1(_2295_),
    .A2(_2299_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5671_ (.A1(_2070_),
    .A2(_2300_),
    .B(_2162_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5672_ (.I(_2131_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5673_ (.A1(_2207_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][3] ),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5674_ (.I(_1904_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5675_ (.A1(_2304_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][3] ),
    .B(_2254_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5676_ (.A1(_2085_),
    .A2(_2130_),
    .B1(_2303_),
    .B2(_2305_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5677_ (.A1(_2302_),
    .A2(_2306_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5678_ (.A1(_2301_),
    .A2(_2307_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5679_ (.I(_2210_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5680_ (.I(_1693_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5681_ (.A1(_2309_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][4] ),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5682_ (.I(_2084_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5683_ (.A1(_2169_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][4] ),
    .B(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5684_ (.A1(_2308_),
    .A2(_2135_),
    .B1(_2310_),
    .B2(_2312_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5685_ (.A1(_2128_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][4] ),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5686_ (.I(_1649_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5687_ (.A1(_2315_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][4] ),
    .B(_2280_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5688_ (.A1(_2277_),
    .A2(_2138_),
    .B1(_2314_),
    .B2(_2316_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5689_ (.A1(_2077_),
    .A2(_2313_),
    .B1(_2317_),
    .B2(_2302_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5690_ (.I(_2318_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5691_ (.A1(_2289_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][5] ),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5692_ (.I(_1768_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5693_ (.A1(_2320_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][5] ),
    .B(_2254_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5694_ (.A1(_2115_),
    .A2(_2141_),
    .A3(_2143_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5695_ (.A1(_2319_),
    .A2(_2321_),
    .B(_2322_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5696_ (.A1(_2095_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][5] ),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5697_ (.I(_1747_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5698_ (.A1(_2325_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][5] ),
    .B(_2084_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5699_ (.A1(_2277_),
    .A2(_2140_),
    .B1(_2324_),
    .B2(_2326_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5700_ (.A1(_2077_),
    .A2(_2323_),
    .B1(_2327_),
    .B2(_2302_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5701_ (.I(_2328_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5702_ (.A1(_2309_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][6] ),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5703_ (.A1(_2169_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][6] ),
    .B(_2311_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5704_ (.A1(_2065_),
    .A2(_2146_),
    .B1(_2329_),
    .B2(_2330_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5705_ (.A1(_2128_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][6] ),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5706_ (.A1(_2315_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][6] ),
    .B(_2280_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5707_ (.A1(_2277_),
    .A2(_2148_),
    .B1(_2332_),
    .B2(_2333_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5708_ (.A1(_2077_),
    .A2(_2331_),
    .B1(_2334_),
    .B2(_2302_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5709_ (.I(_2335_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5710_ (.A1(_2309_),
    .A2(\mod.Data_Mem.F_M.MRAM[29][7] ),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5711_ (.I(_1639_),
    .Z(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5712_ (.I(_2337_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5713_ (.A1(_2338_),
    .A2(\mod.Data_Mem.F_M.MRAM[28][7] ),
    .B(_2311_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5714_ (.A1(_2308_),
    .A2(_2150_),
    .B1(_2336_),
    .B2(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5715_ (.A1(_2278_),
    .A2(\mod.Data_Mem.F_M.MRAM[797][7] ),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5716_ (.A1(_2157_),
    .A2(\mod.Data_Mem.F_M.MRAM[796][7] ),
    .B(_2210_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5717_ (.A1(_2311_),
    .A2(_2152_),
    .B1(_2341_),
    .B2(_2342_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5718_ (.A1(_2062_),
    .A2(_2340_),
    .B1(_2343_),
    .B2(_2164_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5719_ (.I(_2344_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5720_ (.I(_2202_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5721_ (.I(_2345_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5722_ (.A1(_2114_),
    .A2(_1534_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5723_ (.I(_2347_),
    .Z(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5724_ (.A1(_2166_),
    .A2(_1500_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5725_ (.I(_2349_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5726_ (.I(_1695_),
    .Z(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5727_ (.I0(\mod.Data_Mem.F_M.MRAM[14][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][0] ),
    .S(_2351_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5728_ (.I(_1512_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5729_ (.I0(\mod.Data_Mem.F_M.MRAM[16][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][0] ),
    .S(_2353_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5730_ (.I(_2158_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5731_ (.A1(_2110_),
    .A2(_2348_),
    .B1(_2350_),
    .B2(_2352_),
    .C1(_2354_),
    .C2(_2355_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5732_ (.I0(\mod.Data_Mem.F_M.MRAM[4][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[5][0] ),
    .I2(\mod.Data_Mem.F_M.MRAM[20][0] ),
    .I3(\mod.Data_Mem.F_M.MRAM[21][0] ),
    .S0(_1717_),
    .S1(_1757_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5733_ (.I0(\mod.Data_Mem.F_M.MRAM[18][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][0] ),
    .S(_2297_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5734_ (.I(_2058_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5735_ (.I(_2349_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5736_ (.I0(\mod.Data_Mem.F_M.MRAM[2][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][0] ),
    .S(_1971_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5737_ (.A1(_2360_),
    .A2(_2361_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5738_ (.A1(_2359_),
    .A2(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5739_ (.A1(_2355_),
    .A2(_2357_),
    .B1(_2358_),
    .B2(_2348_),
    .C(_2363_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5740_ (.A1(_2346_),
    .A2(_2356_),
    .B(_2364_),
    .C(_1499_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5741_ (.A1(_1547_),
    .A2(_1532_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5742_ (.I(_2366_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5743_ (.A1(_1594_),
    .A2(_1501_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5744_ (.I(_2368_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5745_ (.A1(_2104_),
    .A2(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5746_ (.I(_2370_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5747_ (.I(_2371_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5748_ (.A1(_2087_),
    .A2(_2058_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5749_ (.I(_2373_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5750_ (.I(_2374_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5751_ (.I(_1944_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5752_ (.I0(\mod.Data_Mem.F_M.MRAM[782][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[783][0] ),
    .S(_2376_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5753_ (.I(_2142_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5754_ (.A1(_1717_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][0] ),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5755_ (.A1(_2378_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][0] ),
    .B(_2379_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5756_ (.I(_2099_),
    .Z(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5757_ (.I0(\mod.Data_Mem.F_M.MRAM[770][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][0] ),
    .S(_1915_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5758_ (.I0(\mod.Data_Mem.F_M.MRAM[772][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[773][0] ),
    .S(_1515_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5759_ (.A1(_2381_),
    .A2(_2382_),
    .B1(_2383_),
    .B2(_2273_),
    .C(_2369_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5760_ (.A1(_2203_),
    .A2(_2380_),
    .B(_2384_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5761_ (.A1(_2375_),
    .A2(_2377_),
    .B(_2385_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5762_ (.I(_2373_),
    .Z(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5763_ (.A1(_1594_),
    .A2(_1495_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5764_ (.I(_2388_),
    .Z(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5765_ (.I(_2389_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5766_ (.I(_1840_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5767_ (.A1(_1774_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][0] ),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5768_ (.A1(_2391_),
    .A2(\mod.Data_Mem.F_M.MRAM[788][0] ),
    .B(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5769_ (.A1(_2387_),
    .A2(_2097_),
    .B1(_2390_),
    .B2(_2393_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5770_ (.A1(_2087_),
    .A2(_1553_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5771_ (.I(_2395_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5772_ (.I0(\mod.Data_Mem.F_M.MRAM[784][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][0] ),
    .S(_1956_),
    .Z(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5773_ (.A1(_2396_),
    .A2(_2397_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5774_ (.I(_2107_),
    .Z(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5775_ (.I(_1584_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5776_ (.I0(\mod.Data_Mem.F_M.MRAM[786][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[787][0] ),
    .S(_2400_),
    .Z(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5777_ (.A1(_2399_),
    .A2(_2401_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5778_ (.A1(_2398_),
    .A2(_2402_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5779_ (.A1(_2394_),
    .A2(_2403_),
    .B(_2371_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5780_ (.A1(_2372_),
    .A2(_2386_),
    .B(_2404_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5781_ (.A1(_1490_),
    .A2(_2116_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5782_ (.I(_2406_),
    .Z(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5783_ (.A1(_2073_),
    .A2(_2365_),
    .A3(_2367_),
    .B1(_2405_),
    .B2(_2407_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5784_ (.I(_2408_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5785_ (.I(_2371_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5786_ (.I(_2179_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5787_ (.A1(_2304_),
    .A2(\mod.Data_Mem.F_M.MRAM[787][1] ),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5788_ (.A1(_2410_),
    .A2(_1686_),
    .B(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5789_ (.A1(_2108_),
    .A2(_2412_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5790_ (.I(_1595_),
    .Z(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5791_ (.I(_2414_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5792_ (.A1(_2075_),
    .A2(\mod.Data_Mem.F_M.MRAM[785][1] ),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5793_ (.A1(_2296_),
    .A2(_1683_),
    .B(_2416_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5794_ (.I(_2400_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5795_ (.I(_2388_),
    .Z(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5796_ (.I(_1880_),
    .Z(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5797_ (.A1(_2420_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][1] ),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5798_ (.A1(_2418_),
    .A2(_1689_),
    .B(_2419_),
    .C(_2421_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5799_ (.A1(_2415_),
    .A2(_2121_),
    .B1(_2417_),
    .B2(_2396_),
    .C(_2422_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5800_ (.A1(_2413_),
    .A2(_2423_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5801_ (.I(_1535_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5802_ (.I(_2107_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5803_ (.I(_1835_),
    .Z(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5804_ (.A1(_1791_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][1] ),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5805_ (.A1(_2427_),
    .A2(_1713_),
    .B(_2428_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5806_ (.I0(\mod.Data_Mem.F_M.MRAM[782][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[783][1] ),
    .S(_1711_),
    .Z(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5807_ (.I(_2414_),
    .Z(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5808_ (.I(_2389_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5809_ (.A1(_2209_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][1] ),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5810_ (.I(_2224_),
    .Z(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5811_ (.A1(_2434_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][1] ),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5812_ (.A1(_2432_),
    .A2(_2433_),
    .A3(_2435_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5813_ (.A1(_2426_),
    .A2(_2429_),
    .B1(_2430_),
    .B2(_2431_),
    .C(_2436_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5814_ (.A1(_2425_),
    .A2(_2437_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5815_ (.A1(_2409_),
    .A2(_2424_),
    .B(_2438_),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5816_ (.I(_2088_),
    .Z(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5817_ (.I0(\mod.Data_Mem.F_M.MRAM[4][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[5][1] ),
    .I2(\mod.Data_Mem.F_M.MRAM[20][1] ),
    .I3(\mod.Data_Mem.F_M.MRAM[21][1] ),
    .S0(_1923_),
    .S1(_2104_),
    .Z(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5818_ (.I0(\mod.Data_Mem.F_M.MRAM[2][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][1] ),
    .S(_1786_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5819_ (.I0(\mod.Data_Mem.F_M.MRAM[18][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][1] ),
    .S(_2337_),
    .Z(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5820_ (.I(_2347_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5821_ (.A1(_2440_),
    .A2(_2441_),
    .B1(_2442_),
    .B2(_2360_),
    .C1(_2443_),
    .C2(_2444_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5822_ (.A1(_2346_),
    .A2(_2445_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5823_ (.I(_2359_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5824_ (.I0(\mod.Data_Mem.F_M.MRAM[30][1] ),
    .I1(_1634_),
    .S(_1921_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5825_ (.I0(\mod.Data_Mem.F_M.MRAM[14][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][1] ),
    .S(_1786_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5826_ (.I0(\mod.Data_Mem.F_M.MRAM[16][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][1] ),
    .S(_2337_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5827_ (.A1(_2448_),
    .A2(_2444_),
    .B1(_2350_),
    .B2(_2449_),
    .C1(_2450_),
    .C2(_2168_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5828_ (.A1(_2447_),
    .A2(_2451_),
    .B(_1807_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5829_ (.A1(_2446_),
    .A2(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5830_ (.A1(_2081_),
    .A2(_2439_),
    .B(_2453_),
    .C(_1499_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5831_ (.I(_2107_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5832_ (.A1(_2304_),
    .A2(\mod.Data_Mem.F_M.MRAM[787][2] ),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5833_ (.A1(_2410_),
    .A2(_1793_),
    .B(_2455_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5834_ (.A1(_2454_),
    .A2(_2456_),
    .ZN(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5835_ (.A1(_2325_),
    .A2(\mod.Data_Mem.F_M.MRAM[785][2] ),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5836_ (.A1(_2296_),
    .A2(_1797_),
    .B(_2458_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5837_ (.A1(_2420_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][2] ),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5838_ (.A1(_2418_),
    .A2(_1788_),
    .B(_2419_),
    .C(_2460_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5839_ (.A1(_2431_),
    .A2(_2124_),
    .B1(_2459_),
    .B2(_2396_),
    .C(_2461_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5840_ (.A1(_2457_),
    .A2(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5841_ (.I(_1681_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5842_ (.A1(_2157_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][2] ),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5843_ (.A1(_2464_),
    .A2(_1770_),
    .B(_2465_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5844_ (.I0(\mod.Data_Mem.F_M.MRAM[782][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[783][2] ),
    .S(_1954_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5845_ (.A1(_2209_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][2] ),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5846_ (.A1(_2434_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][2] ),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5847_ (.A1(_2432_),
    .A2(_2468_),
    .A3(_2469_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5848_ (.A1(_2426_),
    .A2(_2466_),
    .B1(_2467_),
    .B2(_2431_),
    .C(_2470_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5849_ (.A1(_2425_),
    .A2(_2471_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5850_ (.A1(_2372_),
    .A2(_2463_),
    .B(_2472_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5851_ (.I0(\mod.Data_Mem.F_M.MRAM[4][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[5][2] ),
    .I2(\mod.Data_Mem.F_M.MRAM[20][2] ),
    .I3(\mod.Data_Mem.F_M.MRAM[21][2] ),
    .S0(_1769_),
    .S1(_2104_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5852_ (.I0(\mod.Data_Mem.F_M.MRAM[2][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][2] ),
    .S(_1786_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5853_ (.I0(\mod.Data_Mem.F_M.MRAM[18][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][2] ),
    .S(_1796_),
    .Z(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5854_ (.A1(_2440_),
    .A2(_2474_),
    .B1(_2475_),
    .B2(_2360_),
    .C1(_2476_),
    .C2(_2444_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5855_ (.A1(_2346_),
    .A2(_2477_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5856_ (.I0(\mod.Data_Mem.F_M.MRAM[14][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][2] ),
    .S(_1774_),
    .Z(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5857_ (.I0(\mod.Data_Mem.F_M.MRAM[16][2] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][2] ),
    .S(_2337_),
    .Z(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5858_ (.A1(_2123_),
    .A2(_2444_),
    .B1(_2360_),
    .B2(_2479_),
    .C1(_2480_),
    .C2(_2168_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5859_ (.A1(_2447_),
    .A2(_2481_),
    .B(_1807_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5860_ (.A1(_2478_),
    .A2(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5861_ (.A1(_2081_),
    .A2(_2473_),
    .B(_2483_),
    .C(_1499_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5862_ (.I(_2381_),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5863_ (.I0(\mod.Data_Mem.F_M.MRAM[786][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[787][3] ),
    .S(_2376_),
    .Z(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5864_ (.A1(_2484_),
    .A2(_2485_),
    .B(_2371_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5865_ (.I(_2388_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5866_ (.I(_2487_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5867_ (.I0(\mod.Data_Mem.F_M.MRAM[788][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[789][3] ),
    .S(_2427_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5868_ (.I(_1712_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5869_ (.I0(\mod.Data_Mem.F_M.MRAM[784][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][3] ),
    .S(_2490_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5870_ (.I(_2369_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5871_ (.A1(_2488_),
    .A2(_2489_),
    .B1(_2491_),
    .B2(_2492_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5872_ (.A1(_2415_),
    .A2(_2130_),
    .B(_2486_),
    .C(_2493_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5873_ (.A1(_2261_),
    .A2(\mod.Data_Mem.F_M.MRAM[782][3] ),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5874_ (.I(_2202_),
    .Z(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5875_ (.A1(_2056_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][3] ),
    .B(_2495_),
    .C(_2496_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5876_ (.I(_2099_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5877_ (.I(_2498_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5878_ (.I(_1791_),
    .Z(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5879_ (.A1(_2296_),
    .A2(\mod.Data_Mem.F_M.MRAM[771][3] ),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5880_ (.A1(_2500_),
    .A2(_1851_),
    .B(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5881_ (.I(_1845_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5882_ (.A1(_2503_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][3] ),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5883_ (.A1(_2338_),
    .A2(_1846_),
    .B(_2504_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5884_ (.I(_2115_),
    .Z(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5885_ (.A1(_2499_),
    .A2(_2502_),
    .B1(_2505_),
    .B2(_2506_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5886_ (.A1(_2372_),
    .A2(_2497_),
    .A3(_2507_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5887_ (.A1(_2117_),
    .A2(_2494_),
    .A3(_2508_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5888_ (.I(_2158_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5889_ (.I0(\mod.Data_Mem.F_M.MRAM[4][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[5][3] ),
    .I2(\mod.Data_Mem.F_M.MRAM[20][3] ),
    .I3(\mod.Data_Mem.F_M.MRAM[21][3] ),
    .S0(_1796_),
    .S1(_1757_),
    .Z(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5890_ (.I0(\mod.Data_Mem.F_M.MRAM[18][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][3] ),
    .S(_2427_),
    .Z(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5891_ (.I0(\mod.Data_Mem.F_M.MRAM[2][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][3] ),
    .S(_2420_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5892_ (.A1(_2510_),
    .A2(_2511_),
    .B1(_2512_),
    .B2(_2348_),
    .C1(_2513_),
    .C2(_2350_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5893_ (.A1(_2204_),
    .A2(_2514_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5894_ (.I(_1944_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5895_ (.I0(\mod.Data_Mem.F_M.MRAM[14][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][3] ),
    .S(_2516_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5896_ (.I0(\mod.Data_Mem.F_M.MRAM[16][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][3] ),
    .S(_2516_),
    .Z(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5897_ (.A1(_2126_),
    .A2(_2348_),
    .B1(_2350_),
    .B2(_2517_),
    .C1(_2518_),
    .C2(_2355_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5898_ (.I(_2116_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5899_ (.A1(_2447_),
    .A2(_2519_),
    .B(_2520_),
    .C(_2219_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5900_ (.A1(_2515_),
    .A2(_2521_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5901_ (.A1(_2074_),
    .A2(_2509_),
    .B(_2522_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5902_ (.I(_1728_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5903_ (.I(_2374_),
    .Z(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5904_ (.I(_2432_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5905_ (.I(_2400_),
    .Z(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5906_ (.A1(_2526_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][4] ),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5907_ (.A1(_2056_),
    .A2(\mod.Data_Mem.F_M.MRAM[788][4] ),
    .B(_2527_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5908_ (.I(_2395_),
    .Z(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5909_ (.I0(\mod.Data_Mem.F_M.MRAM[784][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][4] ),
    .S(_2516_),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5910_ (.A1(_2196_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][4] ),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5911_ (.A1(_2378_),
    .A2(_1922_),
    .B(_2531_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5912_ (.A1(_2529_),
    .A2(_2530_),
    .B1(_2532_),
    .B2(_2426_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5913_ (.A1(_2524_),
    .A2(_2138_),
    .B1(_2525_),
    .B2(_2528_),
    .C(_2533_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5914_ (.I(_2098_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5915_ (.I0(\mod.Data_Mem.F_M.MRAM[782][4] ),
    .I1(_1902_),
    .S(_2434_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5916_ (.I0(\mod.Data_Mem.F_M.MRAM[770][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][4] ),
    .S(_2490_),
    .Z(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5917_ (.I(_2389_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5918_ (.A1(_2259_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][4] ),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5919_ (.I(_1835_),
    .Z(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5920_ (.A1(_2540_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][4] ),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5921_ (.A1(_2538_),
    .A2(_2539_),
    .A3(_2541_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5922_ (.A1(_2415_),
    .A2(_2536_),
    .B1(_2537_),
    .B2(_2454_),
    .C(_2542_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5923_ (.A1(_2535_),
    .A2(_2543_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5924_ (.A1(_2409_),
    .A2(_2534_),
    .B(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5925_ (.I0(\mod.Data_Mem.F_M.MRAM[18][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][4] ),
    .S(_2353_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5926_ (.A1(_2359_),
    .A2(_2546_),
    .B(_2098_),
    .C(_2440_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5927_ (.I(_2395_),
    .Z(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5928_ (.I0(\mod.Data_Mem.F_M.MRAM[16][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][4] ),
    .S(_2353_),
    .Z(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5929_ (.I(_2389_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5930_ (.A1(_2304_),
    .A2(\mod.Data_Mem.F_M.MRAM[21][4] ),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5931_ (.A1(_2269_),
    .A2(\mod.Data_Mem.F_M.MRAM[20][4] ),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5932_ (.A1(_2550_),
    .A2(_2551_),
    .A3(_2552_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5933_ (.A1(_2548_),
    .A2(_2549_),
    .B(_2553_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5934_ (.I(_2059_),
    .Z(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5935_ (.A1(_1532_),
    .A2(_2135_),
    .B1(_2547_),
    .B2(_2554_),
    .C(_2555_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5936_ (.I(_2370_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5937_ (.I(_2434_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5938_ (.I(_2100_),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5939_ (.A1(_2136_),
    .A2(\mod.Data_Mem.F_M.MRAM[3][4] ),
    .Z(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5940_ (.A1(_2558_),
    .A2(\mod.Data_Mem.F_M.MRAM[2][4] ),
    .B(_2559_),
    .C(_2560_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5941_ (.I(_2207_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5942_ (.A1(_2503_),
    .A2(\mod.Data_Mem.F_M.MRAM[4][4] ),
    .Z(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5943_ (.A1(_2562_),
    .A2(\mod.Data_Mem.F_M.MRAM[5][4] ),
    .B(_2563_),
    .C(_2510_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5944_ (.A1(_2503_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][4] ),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5945_ (.A1(_2562_),
    .A2(_1870_),
    .B(_2069_),
    .C(_2565_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5946_ (.A1(_2557_),
    .A2(_2561_),
    .A3(_2564_),
    .A4(_2566_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5947_ (.A1(_2520_),
    .A2(_2556_),
    .A3(_2567_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5948_ (.A1(_2523_),
    .A2(_2545_),
    .B1(_2568_),
    .B2(_2407_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5949_ (.I0(\mod.Data_Mem.F_M.MRAM[18][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[19][5] ),
    .S(_2427_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5950_ (.A1(_2447_),
    .A2(_2569_),
    .B(_1536_),
    .C(_2355_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5951_ (.I(_1712_),
    .Z(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5952_ (.I0(\mod.Data_Mem.F_M.MRAM[16][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][5] ),
    .S(_2571_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5953_ (.A1(_2526_),
    .A2(\mod.Data_Mem.F_M.MRAM[21][5] ),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5954_ (.A1(_2391_),
    .A2(\mod.Data_Mem.F_M.MRAM[20][5] ),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5955_ (.A1(_2390_),
    .A2(_2573_),
    .A3(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5956_ (.A1(_2548_),
    .A2(_2572_),
    .B(_2575_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5957_ (.A1(_1628_),
    .A2(_2141_),
    .A3(_2143_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5958_ (.A1(_2570_),
    .A2(_2576_),
    .B(_2577_),
    .C(_2258_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5959_ (.I(_2269_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5960_ (.A1(_2464_),
    .A2(\mod.Data_Mem.F_M.MRAM[4][5] ),
    .Z(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5961_ (.A1(_2579_),
    .A2(\mod.Data_Mem.F_M.MRAM[5][5] ),
    .B(_2580_),
    .C(_2506_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5962_ (.I(_1512_),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5963_ (.I0(\mod.Data_Mem.F_M.MRAM[2][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][5] ),
    .S(_2582_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5964_ (.I0(\mod.Data_Mem.F_M.MRAM[14][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][5] ),
    .S(_2516_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5965_ (.A1(_2499_),
    .A2(_2583_),
    .B1(_2584_),
    .B2(_2555_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5966_ (.A1(_2557_),
    .A2(_2581_),
    .A3(_2585_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5967_ (.A1(_2520_),
    .A2(_2578_),
    .A3(_2586_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5968_ (.A1(_1774_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][5] ),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5969_ (.A1(_2391_),
    .A2(\mod.Data_Mem.F_M.MRAM[782][5] ),
    .B(_2588_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5970_ (.I(_1840_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5971_ (.A1(_2351_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][5] ),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5972_ (.A1(_2590_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][5] ),
    .B(_2591_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5973_ (.A1(_2387_),
    .A2(_2589_),
    .B1(_2592_),
    .B2(_2390_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5974_ (.I0(\mod.Data_Mem.F_M.MRAM[770][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][5] ),
    .S(_2490_),
    .Z(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5975_ (.A1(_2351_),
    .A2(_1938_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5976_ (.A1(_2540_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][5] ),
    .B(_2595_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5977_ (.I0(\mod.Data_Mem.F_M.MRAM[786][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[787][5] ),
    .S(_1515_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5978_ (.I0(\mod.Data_Mem.F_M.MRAM[784][5] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][5] ),
    .S(_2224_),
    .Z(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5979_ (.A1(_2399_),
    .A2(_2597_),
    .B1(_2598_),
    .B2(_2396_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5980_ (.A1(_2387_),
    .A2(_2140_),
    .B1(_2390_),
    .B2(_2596_),
    .C(_2599_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _5981_ (.A1(_1633_),
    .A2(_2593_),
    .B1(_2594_),
    .B2(_2102_),
    .C1(_2557_),
    .C2(_2600_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5982_ (.A1(_2073_),
    .A2(_2601_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5983_ (.A1(_2407_),
    .A2(_2587_),
    .B(_2602_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5984_ (.I(_2550_),
    .Z(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5985_ (.A1(_2464_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][6] ),
    .Z(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5986_ (.A1(_2579_),
    .A2(\mod.Data_Mem.F_M.MRAM[788][6] ),
    .B(_2604_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5987_ (.A1(_2055_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][6] ),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5988_ (.A1(_2590_),
    .A2(_2009_),
    .B(_2606_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5989_ (.I0(\mod.Data_Mem.F_M.MRAM[784][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][6] ),
    .S(_2297_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5990_ (.A1(_2454_),
    .A2(_2607_),
    .B1(_2608_),
    .B2(_2529_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5991_ (.A1(_2524_),
    .A2(_2148_),
    .B1(_2603_),
    .B2(_2605_),
    .C(_2609_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5992_ (.I(_2136_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5993_ (.A1(_1937_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][6] ),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5994_ (.A1(_2611_),
    .A2(\mod.Data_Mem.F_M.MRAM[782][6] ),
    .B(_2612_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5995_ (.A1(_2418_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][6] ),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5996_ (.A1(_2056_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][6] ),
    .B(_2614_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5997_ (.A1(_2524_),
    .A2(_2613_),
    .B1(_2615_),
    .B2(_2525_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5998_ (.I(_1757_),
    .Z(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5999_ (.I(_2617_),
    .Z(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6000_ (.I0(\mod.Data_Mem.F_M.MRAM[770][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][6] ),
    .S(_2271_),
    .Z(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6001_ (.A1(_2102_),
    .A2(_2619_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6002_ (.A1(_2406_),
    .A2(_2620_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6003_ (.A1(_2409_),
    .A2(_2610_),
    .B1(_2616_),
    .B2(_2618_),
    .C(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6004_ (.I0(\mod.Data_Mem.F_M.MRAM[16][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][6] ),
    .S(_1937_),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6005_ (.A1(_2259_),
    .A2(\mod.Data_Mem.F_M.MRAM[20][6] ),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6006_ (.A1(_2540_),
    .A2(\mod.Data_Mem.F_M.MRAM[21][6] ),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6007_ (.A1(_2538_),
    .A2(_2624_),
    .A3(_2625_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6008_ (.A1(_2400_),
    .A2(\mod.Data_Mem.F_M.MRAM[19][6] ),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6009_ (.A1(_2055_),
    .A2(\mod.Data_Mem.F_M.MRAM[18][6] ),
    .B(_2627_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6010_ (.A1(_2345_),
    .A2(_2628_),
    .B(_2347_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6011_ (.A1(_2548_),
    .A2(_2623_),
    .B(_2626_),
    .C(_2629_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6012_ (.A1(_2183_),
    .A2(_2146_),
    .B(_2630_),
    .C(_2258_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6013_ (.I(_1763_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6014_ (.A1(_2632_),
    .A2(\mod.Data_Mem.F_M.MRAM[4][6] ),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6015_ (.A1(_2579_),
    .A2(\mod.Data_Mem.F_M.MRAM[5][6] ),
    .B(_2633_),
    .C(_2089_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6016_ (.I(_2498_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6017_ (.I0(\mod.Data_Mem.F_M.MRAM[2][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][6] ),
    .S(_2075_),
    .Z(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6018_ (.I0(\mod.Data_Mem.F_M.MRAM[14][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][6] ),
    .S(_2582_),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6019_ (.A1(_2635_),
    .A2(_2636_),
    .B1(_2637_),
    .B2(_2555_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6020_ (.A1(_2372_),
    .A2(_2634_),
    .A3(_2638_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6021_ (.A1(_1676_),
    .A2(_2117_),
    .A3(_2631_),
    .A4(_2639_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6022_ (.A1(_2622_),
    .A2(_2640_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6023_ (.I(_2196_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6024_ (.A1(_2526_),
    .A2(\mod.Data_Mem.F_M.MRAM[789][7] ),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6025_ (.A1(_2641_),
    .A2(\mod.Data_Mem.F_M.MRAM[788][7] ),
    .B(_2642_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6026_ (.I0(\mod.Data_Mem.F_M.MRAM[784][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[785][7] ),
    .S(_2297_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6027_ (.A1(_2196_),
    .A2(\mod.Data_Mem.F_M.MRAM[786][7] ),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6028_ (.A1(_2378_),
    .A2(_2043_),
    .B(_2645_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6029_ (.A1(_2529_),
    .A2(_2644_),
    .B1(_2646_),
    .B2(_2426_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6030_ (.A1(_2524_),
    .A2(_2152_),
    .B1(_2525_),
    .B2(_2643_),
    .C(_2647_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6031_ (.I0(\mod.Data_Mem.F_M.MRAM[782][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[783][7] ),
    .S(_2571_),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6032_ (.I0(\mod.Data_Mem.F_M.MRAM[770][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[771][7] ),
    .S(_2490_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6033_ (.A1(_2540_),
    .A2(\mod.Data_Mem.F_M.MRAM[773][7] ),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6034_ (.A1(_2378_),
    .A2(\mod.Data_Mem.F_M.MRAM[772][7] ),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6035_ (.A1(_2538_),
    .A2(_2651_),
    .A3(_2652_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6036_ (.A1(_2415_),
    .A2(_2649_),
    .B1(_2650_),
    .B2(_2454_),
    .C(_2653_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6037_ (.A1(_2535_),
    .A2(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6038_ (.A1(_2409_),
    .A2(_2648_),
    .B(_2655_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6039_ (.I0(\mod.Data_Mem.F_M.MRAM[16][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[17][7] ),
    .S(_2420_),
    .Z(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6040_ (.A1(_2320_),
    .A2(\mod.Data_Mem.F_M.MRAM[21][7] ),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6041_ (.A1(_2289_),
    .A2(\mod.Data_Mem.F_M.MRAM[20][7] ),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6042_ (.A1(_2432_),
    .A2(_2658_),
    .A3(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6043_ (.A1(_1792_),
    .A2(\mod.Data_Mem.F_M.MRAM[19][7] ),
    .Z(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6044_ (.A1(_2278_),
    .A2(\mod.Data_Mem.F_M.MRAM[18][7] ),
    .B(_2661_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6045_ (.A1(_2345_),
    .A2(_2662_),
    .B(_2347_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6046_ (.A1(_2529_),
    .A2(_2657_),
    .B(_2660_),
    .C(_2663_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6047_ (.A1(_2183_),
    .A2(_2150_),
    .B(_2664_),
    .C(_2258_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6048_ (.I0(\mod.Data_Mem.F_M.MRAM[2][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[3][7] ),
    .S(_2179_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6049_ (.A1(_2635_),
    .A2(_2666_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6050_ (.A1(_2503_),
    .A2(\mod.Data_Mem.F_M.MRAM[4][7] ),
    .Z(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6051_ (.A1(_2562_),
    .A2(\mod.Data_Mem.F_M.MRAM[5][7] ),
    .B(_2668_),
    .C(_2510_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6052_ (.I0(\mod.Data_Mem.F_M.MRAM[14][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[15][7] ),
    .S(_2320_),
    .Z(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6053_ (.A1(_2555_),
    .A2(_2670_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6054_ (.A1(_2557_),
    .A2(_2667_),
    .A3(_2669_),
    .A4(_2671_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6055_ (.A1(_2520_),
    .A2(_2665_),
    .A3(_2672_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6056_ (.A1(_2523_),
    .A2(_2656_),
    .B1(_2673_),
    .B2(_2407_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6057_ (.A1(_1693_),
    .A2(_2395_),
    .B(_1535_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6058_ (.I(_2674_),
    .Z(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6059_ (.A1(_2506_),
    .A2(\mod.Data_Mem.F_M.MRAM[782][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[783][0] ),
    .B2(_2558_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6060_ (.A1(_2675_),
    .A2(_2676_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6061_ (.A1(_1710_),
    .A2(_2368_),
    .B(_1496_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6062_ (.I(_2678_),
    .Z(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6063_ (.I(_2679_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6064_ (.A1(_2170_),
    .A2(_2680_),
    .B(_1731_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6065_ (.I(_2674_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6066_ (.A1(\mod.Data_Mem.F_M.MRAM[797][0] ),
    .A2(_2682_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6067_ (.I(_2678_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6068_ (.I(_2684_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6069_ (.A1(\mod.Data_Mem.F_M.MRAM[781][0] ),
    .A2(_2685_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6070_ (.A1(_2083_),
    .A2(_2683_),
    .A3(_2686_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6071_ (.A1(_2677_),
    .A2(_2681_),
    .B(_1728_),
    .C(_2687_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6072_ (.I(_2271_),
    .Z(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6073_ (.A1(_2689_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[15][0] ),
    .B2(_2506_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6074_ (.A1(\mod.Data_Mem.F_M.MRAM[13][0] ),
    .A2(_2083_),
    .B1(_2205_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][0] ),
    .C(_2105_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6075_ (.A1(_1805_),
    .A2(_2690_),
    .B(_2691_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6076_ (.I(_2079_),
    .Z(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6077_ (.A1(_2076_),
    .A2(_1498_),
    .B1(_2161_),
    .B2(_1633_),
    .C(_2693_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6078_ (.A1(_2202_),
    .A2(_2194_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6079_ (.I(_2695_),
    .Z(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6080_ (.A1(_2692_),
    .A2(_2694_),
    .B(_2696_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6081_ (.I(_1588_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6082_ (.A1(_2698_),
    .A2(_1612_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6083_ (.A1(_1552_),
    .A2(_1546_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6084_ (.I(_2700_),
    .Z(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6085_ (.I(_2701_),
    .Z(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6086_ (.A1(_1830_),
    .A2(_1616_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6087_ (.A1(_2699_),
    .A2(_2702_),
    .A3(_2703_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6088_ (.I(_1873_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6089_ (.A1(_2705_),
    .A2(\mod.Data_Mem.F_M.MRAM[790][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[791][0] ),
    .B2(_2115_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6090_ (.A1(_1648_),
    .A2(_1605_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6091_ (.A1(_1501_),
    .A2(_1545_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6092_ (.I(_2708_),
    .Z(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6093_ (.I(_2709_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6094_ (.A1(_2189_),
    .A2(_2706_),
    .B(_2707_),
    .C(_2710_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6095_ (.A1(_2704_),
    .A2(_2682_),
    .A3(_2711_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6096_ (.I(_2701_),
    .Z(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6097_ (.A1(_2008_),
    .A2(_1586_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6098_ (.A1(_1830_),
    .A2(_1590_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6099_ (.A1(_2713_),
    .A2(_2714_),
    .A3(_2715_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6100_ (.A1(_2705_),
    .A2(\mod.Data_Mem.F_M.MRAM[774][0] ),
    .B1(\mod.Data_Mem.F_M.MRAM[775][0] ),
    .B2(_2158_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6101_ (.A1(_1740_),
    .A2(_1571_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6102_ (.A1(_2177_),
    .A2(_2717_),
    .B(_2718_),
    .C(_2710_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6103_ (.A1(_2685_),
    .A2(_2716_),
    .A3(_2719_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6104_ (.A1(_2183_),
    .A2(_2712_),
    .A3(_2720_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6105_ (.I(_1783_),
    .Z(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6106_ (.A1(_2571_),
    .A2(\mod.Data_Mem.F_M.MRAM[2][0] ),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6107_ (.A1(_2722_),
    .A2(\mod.Data_Mem.F_M.MRAM[3][0] ),
    .B(_1808_),
    .C(_2723_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6108_ (.A1(\mod.Data_Mem.F_M.MRAM[1][0] ),
    .A2(_1539_),
    .B1(_1813_),
    .B2(\mod.Data_Mem.F_M.MRAM[0][0] ),
    .C(_2702_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6109_ (.I0(\mod.Data_Mem.F_M.MRAM[7][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[6][0] ),
    .S(_2179_),
    .Z(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6110_ (.I(_2709_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6111_ (.A1(_1544_),
    .A2(_1506_),
    .B1(_1577_),
    .B2(_2726_),
    .C(_2727_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6112_ (.A1(_2366_),
    .A2(_2680_),
    .B1(_2724_),
    .B2(_2725_),
    .C(_2728_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6113_ (.I0(\mod.Data_Mem.F_M.MRAM[23][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[22][0] ),
    .S(_1717_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6114_ (.A1(_1506_),
    .A2(_1513_),
    .B1(_2730_),
    .B2(_1936_),
    .C(_2727_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6115_ (.A1(_2366_),
    .A2(_2684_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6116_ (.I(_2700_),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6117_ (.A1(_1540_),
    .A2(_1516_),
    .B1(_1520_),
    .B2(_1614_),
    .C(_2733_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6118_ (.A1(_2732_),
    .A2(_2734_),
    .Z(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6119_ (.A1(_2689_),
    .A2(_1498_),
    .B1(_2731_),
    .B2(_2735_),
    .C(_1865_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6120_ (.A1(_2359_),
    .A2(_2189_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6121_ (.A1(_1728_),
    .A2(_2721_),
    .B1(_2729_),
    .B2(_2736_),
    .C(_2737_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6122_ (.A1(_2688_),
    .A2(_2697_),
    .B(_2738_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6123_ (.A1(_2611_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][1] ),
    .B2(_2085_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6124_ (.A1(\mod.Data_Mem.F_M.MRAM[781][1] ),
    .A2(_2193_),
    .B1(_2195_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][1] ),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6125_ (.A1(_2165_),
    .A2(_2739_),
    .B(_2740_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6126_ (.A1(_2182_),
    .A2(_2682_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6127_ (.A1(_2675_),
    .A2(_2741_),
    .B(_2742_),
    .C(_2080_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6128_ (.I(_2684_),
    .Z(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6129_ (.I(_1537_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6130_ (.I(_1525_),
    .Z(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6131_ (.A1(_2114_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[15][1] ),
    .B2(_1944_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6132_ (.A1(_2746_),
    .A2(_2747_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6133_ (.A1(\mod.Data_Mem.F_M.MRAM[13][1] ),
    .A2(_2745_),
    .B1(_2153_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][1] ),
    .C(_2748_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6134_ (.A1(_2744_),
    .A2(_2749_),
    .Z(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6135_ (.A1(_2186_),
    .A2(_2682_),
    .B(_2750_),
    .C(_1865_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6136_ (.A1(_2696_),
    .A2(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6137_ (.I(_2225_),
    .Z(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6138_ (.A1(_2325_),
    .A2(\mod.Data_Mem.F_M.MRAM[6][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[7][1] ),
    .B2(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6139_ (.A1(_1804_),
    .A2(_1640_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6140_ (.A1(_2177_),
    .A2(_2754_),
    .B(_2755_),
    .C(_2710_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6141_ (.I(_2700_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6142_ (.A1(_1602_),
    .A2(_1650_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6143_ (.A1(_1740_),
    .A2(_1652_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6144_ (.A1(_2757_),
    .A2(_2758_),
    .A3(_2759_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6145_ (.A1(_2744_),
    .A2(_2756_),
    .A3(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6146_ (.A1(_1752_),
    .A2(_1663_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6147_ (.A1(_2178_),
    .A2(_1659_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6148_ (.A1(_2757_),
    .A2(_2762_),
    .A3(_2763_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6149_ (.A1(_2582_),
    .A2(\mod.Data_Mem.F_M.MRAM[22][1] ),
    .B1(\mod.Data_Mem.F_M.MRAM[23][1] ),
    .B2(_2753_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6150_ (.A1(_1911_),
    .A2(_1668_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6151_ (.I(_2708_),
    .Z(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6152_ (.A1(_1643_),
    .A2(_2765_),
    .B(_2766_),
    .C(_2767_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6153_ (.A1(_2674_),
    .A2(_2764_),
    .A3(_2768_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6154_ (.A1(_2761_),
    .A2(_2769_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6155_ (.I(_2701_),
    .Z(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6156_ (.I(_1568_),
    .Z(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6157_ (.A1(_1558_),
    .A2(_1705_),
    .B1(_1707_),
    .B2(_2772_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6158_ (.I(_1607_),
    .Z(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6159_ (.A1(_2774_),
    .A2(_1721_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6160_ (.A1(_1733_),
    .A2(_1715_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6161_ (.A1(_2702_),
    .A2(_2775_),
    .A3(_2776_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6162_ (.A1(_2771_),
    .A2(_2773_),
    .B(_2777_),
    .C(_2685_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6163_ (.A1(_1920_),
    .A2(_1697_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6164_ (.A1(_1608_),
    .A2(_1691_),
    .B(_2733_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6165_ (.A1(_2774_),
    .A2(_1685_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6166_ (.I(_2708_),
    .Z(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6167_ (.A1(_1737_),
    .A2(_1688_),
    .B(_2782_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6168_ (.I(_2678_),
    .Z(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6169_ (.A1(_2779_),
    .A2(_2780_),
    .B1(_2781_),
    .B2(_2783_),
    .C(_2784_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6170_ (.A1(_1807_),
    .A2(_2785_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6171_ (.A1(_2219_),
    .A2(_2770_),
    .B1(_2778_),
    .B2(_2786_),
    .C(_2737_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6172_ (.A1(_2743_),
    .A2(_2752_),
    .B(_2787_),
    .C(_2367_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6173_ (.A1(_2192_),
    .A2(_2675_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6174_ (.A1(_2209_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][2] ),
    .B2(_2280_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6175_ (.A1(_2772_),
    .A2(_2789_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6176_ (.A1(\mod.Data_Mem.F_M.MRAM[781][2] ),
    .A2(_1731_),
    .B1(_2195_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][2] ),
    .C(_2790_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6177_ (.A1(_2680_),
    .A2(_2791_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6178_ (.A1(_2067_),
    .A2(_2788_),
    .A3(_2792_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6179_ (.A1(_2199_),
    .A2(_2675_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6180_ (.A1(_2064_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[15][2] ),
    .B2(_2095_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6181_ (.A1(_1589_),
    .A2(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6182_ (.A1(\mod.Data_Mem.F_M.MRAM[13][2] ),
    .A2(_2193_),
    .B1(_1813_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][2] ),
    .C(_2796_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6183_ (.A1(_2680_),
    .A2(_2797_),
    .B(_2693_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6184_ (.A1(_2794_),
    .A2(_2798_),
    .B(_2696_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6185_ (.A1(_2325_),
    .A2(\mod.Data_Mem.F_M.MRAM[6][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[7][2] ),
    .B2(_2753_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6186_ (.A1(_1804_),
    .A2(_1734_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6187_ (.A1(_2177_),
    .A2(_2800_),
    .B(_2801_),
    .C(_2710_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6188_ (.A1(_1752_),
    .A2(_1741_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6189_ (.A1(_2178_),
    .A2(_1738_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6190_ (.A1(_2757_),
    .A2(_2803_),
    .A3(_2804_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6191_ (.A1(_2744_),
    .A2(_2802_),
    .A3(_2805_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6192_ (.A1(_1752_),
    .A2(_1748_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6193_ (.A1(_2178_),
    .A2(_1744_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6194_ (.A1(_2757_),
    .A2(_2807_),
    .A3(_2808_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6195_ (.A1(_2582_),
    .A2(\mod.Data_Mem.F_M.MRAM[22][2] ),
    .B1(\mod.Data_Mem.F_M.MRAM[23][2] ),
    .B2(_2753_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6196_ (.A1(_1882_),
    .A2(_1753_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6197_ (.A1(_1643_),
    .A2(_2810_),
    .B(_2811_),
    .C(_2767_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6198_ (.A1(_2674_),
    .A2(_2809_),
    .A3(_2812_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6199_ (.A1(_2806_),
    .A2(_2813_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6200_ (.A1(_2772_),
    .A2(_1764_),
    .B1(_1765_),
    .B2(_1558_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6201_ (.A1(_2774_),
    .A2(_1777_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6202_ (.A1(_1733_),
    .A2(_1772_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6203_ (.A1(_2702_),
    .A2(_2816_),
    .A3(_2817_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6204_ (.A1(_2771_),
    .A2(_2815_),
    .B(_2818_),
    .C(_2685_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6205_ (.A1(_1920_),
    .A2(_1785_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6206_ (.A1(_1608_),
    .A2(_1790_),
    .B(_2733_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6207_ (.A1(_2774_),
    .A2(_1799_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6208_ (.A1(_1737_),
    .A2(_1795_),
    .B(_2782_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6209_ (.A1(_2820_),
    .A2(_2821_),
    .B1(_2822_),
    .B2(_2823_),
    .C(_2679_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6210_ (.A1(_1899_),
    .A2(_2824_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6211_ (.A1(_2219_),
    .A2(_2814_),
    .B1(_2819_),
    .B2(_2825_),
    .C(_2737_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6212_ (.A1(_2793_),
    .A2(_2799_),
    .B(_2826_),
    .C(_2367_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6213_ (.I(_2105_),
    .Z(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6214_ (.A1(_2205_),
    .A2(_2212_),
    .B(_2496_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6215_ (.A1(_2558_),
    .A2(_2510_),
    .A3(\mod.Data_Mem.F_M.MRAM[20][3] ),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6216_ (.A1(_2828_),
    .A2(_2829_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6217_ (.I0(\mod.Data_Mem.F_M.MRAM[1][3] ),
    .I1(\mod.Data_Mem.F_M.MRAM[2][3] ),
    .I2(\mod.Data_Mem.F_M.MRAM[3][3] ),
    .I3(\mod.Data_Mem.F_M.MRAM[4][3] ),
    .S0(_2632_),
    .S1(_2440_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6218_ (.A1(_1614_),
    .A2(_1820_),
    .Z(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6219_ (.A1(_2709_),
    .A2(_2678_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6220_ (.A1(_1936_),
    .A2(_1818_),
    .B(_2832_),
    .C(_2833_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6221_ (.A1(_2210_),
    .A2(\mod.Data_Mem.F_M.MRAM[14][3] ),
    .B1(\mod.Data_Mem.F_M.MRAM[15][3] ),
    .B2(_2278_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6222_ (.A1(_1569_),
    .A2(_2835_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6223_ (.A1(_1622_),
    .A2(_2695_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6224_ (.A1(\mod.Data_Mem.F_M.MRAM[13][3] ),
    .A2(_2193_),
    .B(_2836_),
    .C(_2837_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6225_ (.A1(_2834_),
    .A2(_2838_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6226_ (.A1(_2827_),
    .A2(_2830_),
    .B1(_2831_),
    .B2(_2091_),
    .C(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6227_ (.A1(_2165_),
    .A2(_1836_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6228_ (.I(_2709_),
    .Z(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6229_ (.A1(_1805_),
    .A2(_1832_),
    .B(_2842_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6230_ (.A1(_1740_),
    .A2(_1828_),
    .Z(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6231_ (.A1(_2156_),
    .A2(_1826_),
    .B(_2771_),
    .C(_2844_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6232_ (.A1(_2841_),
    .A2(_2843_),
    .B(_2732_),
    .C(_2845_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(_1936_),
    .A2(_1848_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6234_ (.A1(_2156_),
    .A2(_1842_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6235_ (.A1(_2842_),
    .A2(_2847_),
    .A3(_2848_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6236_ (.A1(_2156_),
    .A2(_1853_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6237_ (.A1(_1577_),
    .A2(_1857_),
    .B(_2727_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6238_ (.A1(_2850_),
    .A2(_2851_),
    .B(_2732_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6239_ (.A1(_2849_),
    .A2(_2852_),
    .B(_2737_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6240_ (.I(\mod.Data_Mem.F_M.MRAM[781][3] ),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6241_ (.I(_1637_),
    .Z(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6242_ (.A1(_2128_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][3] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][3] ),
    .B2(_2064_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6243_ (.A1(_2854_),
    .A2(_2214_),
    .B1(_2855_),
    .B2(_2856_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6244_ (.A1(_2617_),
    .A2(_2857_),
    .B(_2195_),
    .C(_2203_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6245_ (.A1(_2106_),
    .A2(_2217_),
    .B(_2858_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6246_ (.A1(_2846_),
    .A2(_2853_),
    .B(_2859_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6247_ (.I(_1865_),
    .Z(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6248_ (.A1(_2205_),
    .A2(_1628_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6249_ (.A1(_2861_),
    .A2(_2862_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6250_ (.A1(_2523_),
    .A2(_2840_),
    .B1(_2860_),
    .B2(_2863_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6251_ (.I(_2367_),
    .Z(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6252_ (.I(_2695_),
    .Z(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6253_ (.I(_2865_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6254_ (.I(_2679_),
    .Z(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6255_ (.I(_1581_),
    .Z(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6256_ (.A1(_2868_),
    .A2(_1875_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6257_ (.I(_2700_),
    .Z(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6258_ (.A1(_2698_),
    .A2(_1877_),
    .B(_2870_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6259_ (.A1(_2855_),
    .A2(_1881_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6260_ (.I(_1661_),
    .Z(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6261_ (.A1(_2873_),
    .A2(_1879_),
    .B(_2767_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6262_ (.A1(_2869_),
    .A2(_2871_),
    .B1(_2872_),
    .B2(_2874_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6263_ (.A1(_2867_),
    .A2(_2875_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6264_ (.I0(_1891_),
    .I1(_1893_),
    .S(_1746_),
    .Z(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6265_ (.A1(_2701_),
    .A2(_2684_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6266_ (.I(_2878_),
    .Z(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6267_ (.I0(_1895_),
    .I1(_1894_),
    .S(_1896_),
    .Z(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6268_ (.I(_2833_),
    .Z(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6269_ (.A1(_2877_),
    .A2(_2879_),
    .B1(_2880_),
    .B2(_2881_),
    .C(_2072_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6270_ (.I(_2679_),
    .Z(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6271_ (.A1(_2868_),
    .A2(_1905_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6272_ (.A1(_1638_),
    .A2(_1907_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6273_ (.A1(_2842_),
    .A2(_2884_),
    .A3(_2885_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6274_ (.I(_1637_),
    .Z(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6275_ (.A1(_2887_),
    .A2(_1910_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6276_ (.I(_1581_),
    .Z(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6277_ (.A1(_2889_),
    .A2(_1909_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6278_ (.A1(_2713_),
    .A2(_2888_),
    .A3(_2890_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6279_ (.A1(_2883_),
    .A2(_2886_),
    .A3(_2891_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6280_ (.I(_2878_),
    .Z(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6281_ (.I0(\mod.Data_Mem.F_M.MRAM[789][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[791][4] ),
    .I2(\mod.Data_Mem.F_M.MRAM[790][4] ),
    .I3(\mod.Data_Mem.F_M.MRAM[788][4] ),
    .S0(_2167_),
    .S1(_2376_),
    .Z(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6282_ (.I(_1607_),
    .Z(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6283_ (.I0(_1925_),
    .I1(_1926_),
    .S(_2895_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6284_ (.I(_2833_),
    .Z(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6285_ (.A1(_2893_),
    .A2(_2894_),
    .B1(_2896_),
    .B2(_2897_),
    .C(_1899_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6286_ (.A1(_2876_),
    .A2(_2882_),
    .B1(_2892_),
    .B2(_2898_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6287_ (.I(_1537_),
    .Z(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6288_ (.I(_1546_),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6289_ (.I(_1525_),
    .Z(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6290_ (.I(_2053_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6291_ (.I(_1493_),
    .Z(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6292_ (.A1(_2903_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][4] ),
    .B1(\mod.Data_Mem.F_M.MRAM[14][4] ),
    .B2(_2904_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6293_ (.A1(_2902_),
    .A2(_2905_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6294_ (.A1(\mod.Data_Mem.F_M.MRAM[13][4] ),
    .A2(_2900_),
    .B1(_2901_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][4] ),
    .C(_2906_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6295_ (.A1(_2142_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][4] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][4] ),
    .B2(_1494_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6296_ (.A1(_2746_),
    .A2(_2908_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6297_ (.A1(\mod.Data_Mem.F_M.MRAM[781][4] ),
    .A2(_2745_),
    .B1(_2153_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][4] ),
    .C(_2909_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6298_ (.I0(_2228_),
    .I1(_2232_),
    .I2(_2907_),
    .I3(_2910_),
    .S0(_2079_),
    .S1(_2744_),
    .Z(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6299_ (.A1(_2696_),
    .A2(_2911_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6300_ (.A1(_2866_),
    .A2(_2899_),
    .B(_2912_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6301_ (.A1(_2864_),
    .A2(_2913_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6302_ (.A1(_2868_),
    .A2(_1966_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6303_ (.A1(_2698_),
    .A2(_1967_),
    .B(_2870_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6304_ (.A1(_2855_),
    .A2(_1972_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6305_ (.A1(_2873_),
    .A2(_1970_),
    .B(_2782_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6306_ (.A1(_2914_),
    .A2(_2915_),
    .B1(_2916_),
    .B2(_2917_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6307_ (.A1(_2867_),
    .A2(_2918_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6308_ (.I0(_1976_),
    .I1(_1977_),
    .S(_1746_),
    .Z(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6309_ (.I0(_1978_),
    .I1(_1979_),
    .S(_1839_),
    .Z(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6310_ (.A1(_2893_),
    .A2(_2920_),
    .B1(_2921_),
    .B2(_2881_),
    .C(_2072_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6311_ (.A1(_1577_),
    .A2(_1952_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6312_ (.A1(_1657_),
    .A2(_1953_),
    .B(_2870_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6313_ (.A1(_2923_),
    .A2(_2924_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6314_ (.A1(_1638_),
    .A2(_1959_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6315_ (.A1(_2889_),
    .A2(_1958_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6316_ (.A1(_2713_),
    .A2(_2926_),
    .A3(_2927_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6317_ (.A1(_2883_),
    .A2(_2925_),
    .A3(_2928_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6318_ (.A1(_1737_),
    .A2(_1941_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6319_ (.A1(_2772_),
    .A2(_1940_),
    .B(_2930_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6320_ (.I0(_1945_),
    .I1(_1947_),
    .S(_2895_),
    .Z(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6321_ (.A1(_2879_),
    .A2(_2931_),
    .B1(_2932_),
    .B2(_2897_),
    .C(_1675_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6322_ (.A1(_2919_),
    .A2(_2922_),
    .B1(_2929_),
    .B2(_2933_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6323_ (.A1(_2903_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][5] ),
    .B1(\mod.Data_Mem.F_M.MRAM[14][5] ),
    .B2(_2253_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6324_ (.A1(_2902_),
    .A2(_2935_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6325_ (.A1(\mod.Data_Mem.F_M.MRAM[13][5] ),
    .A2(_2900_),
    .B1(_2901_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][5] ),
    .C(_2936_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6326_ (.A1(_2268_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][5] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][5] ),
    .B2(_2904_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6327_ (.A1(_2746_),
    .A2(_2938_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6328_ (.A1(\mod.Data_Mem.F_M.MRAM[781][5] ),
    .A2(_2745_),
    .B1(_2153_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][5] ),
    .C(_2939_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6329_ (.I0(_2235_),
    .I1(_2238_),
    .I2(_2937_),
    .I3(_2940_),
    .S0(_2079_),
    .S1(_2784_),
    .Z(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6330_ (.A1(_2865_),
    .A2(_2941_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6331_ (.A1(_2866_),
    .A2(_2934_),
    .B(_2942_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6332_ (.A1(_2864_),
    .A2(_2943_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6333_ (.A1(_1582_),
    .A2(_2002_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6334_ (.A1(_2887_),
    .A2(_2003_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6335_ (.A1(_2842_),
    .A2(_2944_),
    .A3(_2945_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6336_ (.A1(_1569_),
    .A2(_2001_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6337_ (.A1(_1582_),
    .A2(_2000_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6338_ (.A1(_2771_),
    .A2(_2947_),
    .A3(_2948_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6339_ (.A1(_2883_),
    .A2(_2946_),
    .A3(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6340_ (.I0(\mod.Data_Mem.F_M.MRAM[789][6] ),
    .I1(\mod.Data_Mem.F_M.MRAM[791][6] ),
    .I2(\mod.Data_Mem.F_M.MRAM[790][6] ),
    .I3(\mod.Data_Mem.F_M.MRAM[788][6] ),
    .S0(_2167_),
    .S1(_2315_),
    .Z(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6341_ (.I0(_2011_),
    .I1(_2012_),
    .S(_1839_),
    .Z(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6342_ (.A1(_2893_),
    .A2(_2951_),
    .B1(_2952_),
    .B2(_2881_),
    .C(_1899_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6343_ (.A1(_2855_),
    .A2(_1988_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6344_ (.A1(_1662_),
    .A2(_1987_),
    .B(_2782_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6345_ (.A1(_2873_),
    .A2(_1985_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6346_ (.A1(_1920_),
    .A2(_1986_),
    .B(_2733_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6347_ (.A1(_2954_),
    .A2(_2955_),
    .B1(_2956_),
    .B2(_2957_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6348_ (.A1(_2867_),
    .A2(_2958_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6349_ (.I0(_1995_),
    .I1(_1994_),
    .S(_1844_),
    .Z(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6350_ (.I0(_1992_),
    .I1(_1993_),
    .S(_2895_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6351_ (.A1(_2881_),
    .A2(_2960_),
    .B1(_2961_),
    .B2(_2879_),
    .C(_1727_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6352_ (.A1(_2950_),
    .A2(_2953_),
    .B1(_2959_),
    .B2(_2962_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6353_ (.A1(_2903_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][6] ),
    .B1(\mod.Data_Mem.F_M.MRAM[14][6] ),
    .B2(_2253_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6354_ (.A1(_2902_),
    .A2(_2964_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6355_ (.A1(\mod.Data_Mem.F_M.MRAM[13][6] ),
    .A2(_2900_),
    .B1(_2194_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][6] ),
    .C(_2965_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6356_ (.A1(_2268_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][6] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][6] ),
    .B2(_2904_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6357_ (.A1(_2746_),
    .A2(_2967_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6358_ (.A1(\mod.Data_Mem.F_M.MRAM[781][6] ),
    .A2(_2745_),
    .B1(_2901_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][6] ),
    .C(_2968_),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6359_ (.I0(_2241_),
    .I1(_2244_),
    .I2(_2966_),
    .I3(_2969_),
    .S0(_1489_),
    .S1(_2784_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6360_ (.A1(_2865_),
    .A2(_2970_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6361_ (.A1(_2866_),
    .A2(_2963_),
    .B(_2971_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6362_ (.A1(_2864_),
    .A2(_2972_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6363_ (.A1(_2887_),
    .A2(_2021_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6364_ (.A1(_2873_),
    .A2(_2020_),
    .B(_2767_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6365_ (.A1(_2889_),
    .A2(_2022_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6366_ (.A1(_2698_),
    .A2(_2023_),
    .B(_2870_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6367_ (.A1(_2973_),
    .A2(_2974_),
    .B1(_2975_),
    .B2(_2976_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6368_ (.A1(_2867_),
    .A2(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6369_ (.I0(_2027_),
    .I1(_2028_),
    .S(_1746_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6370_ (.I0(_2029_),
    .I1(_2030_),
    .S(_2895_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6371_ (.A1(_2893_),
    .A2(_2979_),
    .B1(_2980_),
    .B2(_2897_),
    .C(_2072_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6372_ (.A1(_2887_),
    .A2(_2036_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6373_ (.A1(_2889_),
    .A2(_2035_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6374_ (.A1(_2713_),
    .A2(_2982_),
    .A3(_2983_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6375_ (.A1(_2868_),
    .A2(_2037_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6376_ (.A1(_1638_),
    .A2(_2038_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6377_ (.A1(_2727_),
    .A2(_2985_),
    .A3(_2986_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6378_ (.A1(_2883_),
    .A2(_2984_),
    .A3(_2987_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6379_ (.I0(\mod.Data_Mem.F_M.MRAM[789][7] ),
    .I1(\mod.Data_Mem.F_M.MRAM[791][7] ),
    .I2(\mod.Data_Mem.F_M.MRAM[790][7] ),
    .I3(\mod.Data_Mem.F_M.MRAM[788][7] ),
    .S0(_2167_),
    .S1(_2376_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6380_ (.I0(_2045_),
    .I1(_2046_),
    .S(_1804_),
    .Z(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6381_ (.A1(_2879_),
    .A2(_2989_),
    .B1(_2990_),
    .B2(_2897_),
    .C(_1675_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6382_ (.A1(_2978_),
    .A2(_2981_),
    .B1(_2988_),
    .B2(_2991_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6383_ (.A1(_2903_),
    .A2(\mod.Data_Mem.F_M.MRAM[15][7] ),
    .B1(\mod.Data_Mem.F_M.MRAM[14][7] ),
    .B2(_2253_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6384_ (.A1(_1568_),
    .A2(_2993_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6385_ (.A1(\mod.Data_Mem.F_M.MRAM[13][7] ),
    .A2(_1538_),
    .B1(_2194_),
    .B2(\mod.Data_Mem.F_M.MRAM[12][7] ),
    .C(_2994_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6386_ (.A1(_2268_),
    .A2(\mod.Data_Mem.F_M.MRAM[783][7] ),
    .B1(\mod.Data_Mem.F_M.MRAM[782][7] ),
    .B2(_2904_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6387_ (.A1(_2902_),
    .A2(_2996_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6388_ (.A1(\mod.Data_Mem.F_M.MRAM[781][7] ),
    .A2(_2900_),
    .B1(_2901_),
    .B2(\mod.Data_Mem.F_M.MRAM[780][7] ),
    .C(_2997_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6389_ (.I0(_2247_),
    .I1(_2250_),
    .I2(_2995_),
    .I3(_2998_),
    .S0(_1489_),
    .S1(_2784_),
    .Z(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6390_ (.A1(_2865_),
    .A2(_2999_),
    .ZN(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6391_ (.A1(_2866_),
    .A2(_2992_),
    .B(_3000_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6392_ (.A1(_2864_),
    .A2(_3001_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6393_ (.I(_2617_),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6394_ (.I(_2090_),
    .Z(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6395_ (.I(_2419_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6396_ (.I(_2381_),
    .Z(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6397_ (.A1(_3003_),
    .A2(_2256_),
    .B1(_3004_),
    .B2(_2401_),
    .C1(_2397_),
    .C2(_3005_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6398_ (.A1(_3002_),
    .A2(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6399_ (.I(_2487_),
    .Z(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6400_ (.A1(_2705_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][0] ),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6401_ (.A1(_2207_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][0] ),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6402_ (.A1(_2414_),
    .A2(_3009_),
    .A3(_3010_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6403_ (.A1(_3008_),
    .A2(_2382_),
    .B1(_2377_),
    .B2(_2492_),
    .C(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6404_ (.I(_2098_),
    .Z(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6405_ (.A1(_2108_),
    .A2(_2380_),
    .B(_3012_),
    .C(_3013_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6406_ (.A1(_2861_),
    .A2(_3007_),
    .A3(_3014_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6407_ (.I(_2590_),
    .Z(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6408_ (.A1(_2500_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][0] ),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6409_ (.A1(_3016_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][0] ),
    .B(_2375_),
    .C(_3017_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6410_ (.I(_2369_),
    .Z(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6411_ (.I(_3019_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6412_ (.I0(\mod.Data_Mem.F_M.MRAM[0][0] ),
    .I1(\mod.Data_Mem.F_M.MRAM[1][0] ),
    .S(_2705_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6413_ (.I(_2381_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6414_ (.I(_2487_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6415_ (.A1(_3020_),
    .A2(_2352_),
    .B1(_3021_),
    .B2(_3022_),
    .C1(_3023_),
    .C2(_2361_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6416_ (.A1(_2535_),
    .A2(_3018_),
    .A3(_3024_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6417_ (.I(_2419_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6418_ (.A1(_2346_),
    .A2(_2266_),
    .B1(_2358_),
    .B2(_3026_),
    .C1(_2354_),
    .C2(_2499_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6419_ (.A1(_2618_),
    .A2(_3027_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6420_ (.A1(_1762_),
    .A2(_3025_),
    .A3(_3028_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6421_ (.A1(_3015_),
    .A2(_3029_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6422_ (.I(_2090_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6423_ (.A1(_3030_),
    .A2(_2275_),
    .B1(_3023_),
    .B2(_2412_),
    .C1(_2417_),
    .C2(_3022_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6424_ (.A1(_3019_),
    .A2(_2430_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6425_ (.A1(_2353_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][1] ),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6426_ (.A1(_2309_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][1] ),
    .B(_2374_),
    .C(_3033_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6427_ (.A1(_1767_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][1] ),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6428_ (.A1(_1937_),
    .A2(_1719_),
    .B(_3035_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6429_ (.A1(_2550_),
    .A2(_2429_),
    .B1(_3036_),
    .B2(_2498_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6430_ (.A1(_1536_),
    .A2(_3032_),
    .A3(_3034_),
    .A4(_3037_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6431_ (.A1(_2693_),
    .A2(_3038_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6432_ (.A1(_2618_),
    .A2(_3031_),
    .B(_3039_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6433_ (.A1(_2590_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][1] ),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6434_ (.A1(_2632_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][1] ),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6435_ (.A1(_2065_),
    .A2(_3041_),
    .A3(_3042_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6436_ (.A1(_2308_),
    .A2(_2449_),
    .B(_3043_),
    .C(_3003_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6437_ (.I0(\mod.Data_Mem.F_M.MRAM[0][1] ),
    .I1(\mod.Data_Mem.F_M.MRAM[1][1] ),
    .S(_2252_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6438_ (.A1(_3026_),
    .A2(_2442_),
    .B1(_3045_),
    .B2(_3005_),
    .C(_1623_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6439_ (.I(_2090_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6440_ (.A1(_3047_),
    .A2(_2282_),
    .B1(_3008_),
    .B2(_2443_),
    .C1(_2450_),
    .C2(_2484_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6441_ (.I(_2105_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6442_ (.A1(_3044_),
    .A2(_3046_),
    .B1(_3048_),
    .B2(_3049_),
    .C(_2080_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6443_ (.A1(_3040_),
    .A2(_3050_),
    .Z(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6444_ (.I(_3051_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6445_ (.A1(_3030_),
    .A2(_2287_),
    .B1(_3004_),
    .B2(_2456_),
    .C1(_2459_),
    .C2(_3022_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6446_ (.A1(_3002_),
    .A2(_3052_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6447_ (.A1(_3016_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][2] ),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6448_ (.A1(_2689_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][2] ),
    .B(_2375_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6449_ (.A1(_2320_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][2] ),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6450_ (.A1(_2410_),
    .A2(_1775_),
    .B(_3056_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6451_ (.I(_2100_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6452_ (.I(_2487_),
    .Z(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6453_ (.A1(_2492_),
    .A2(_2467_),
    .B1(_3057_),
    .B2(_3058_),
    .C1(_3059_),
    .C2(_2466_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6454_ (.A1(_3054_),
    .A2(_3055_),
    .B(_3060_),
    .C(_3013_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6455_ (.A1(_2861_),
    .A2(_3053_),
    .A3(_3061_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6456_ (.I(_2498_),
    .Z(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6457_ (.A1(\mod.Data_Mem.F_M.MRAM[13][2] ),
    .A2(_2375_),
    .B1(_3063_),
    .B2(\mod.Data_Mem.F_M.MRAM[1][2] ),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6458_ (.A1(_2057_),
    .A2(_3064_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6459_ (.A1(_2722_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][2] ),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6460_ (.A1(_3020_),
    .A2(_2479_),
    .B1(_3066_),
    .B2(_3063_),
    .C(_1633_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6461_ (.A1(\mod.Data_Mem.F_M.MRAM[12][2] ),
    .A2(_1886_),
    .B1(_2525_),
    .B2(_2475_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6462_ (.A1(_3067_),
    .A2(_3068_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6463_ (.A1(_3047_),
    .A2(_2293_),
    .B1(_3008_),
    .B2(_2476_),
    .C1(_2480_),
    .C2(_2484_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6464_ (.A1(_2827_),
    .A2(_3070_),
    .B(_2080_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6465_ (.A1(_3065_),
    .A2(_3069_),
    .B(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6466_ (.A1(_3062_),
    .A2(_3072_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6467_ (.A1(_2169_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][3] ),
    .Z(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6468_ (.A1(_3016_),
    .A2(\mod.Data_Mem.F_M.MRAM[1][3] ),
    .B(_2635_),
    .C(_3073_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6469_ (.A1(_2259_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][3] ),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6470_ (.A1(_2261_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][3] ),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6471_ (.A1(_2414_),
    .A2(_3075_),
    .A3(_3076_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6472_ (.A1(_3020_),
    .A2(_2517_),
    .B1(_2513_),
    .B2(_3004_),
    .C(_3077_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6473_ (.A1(_2535_),
    .A2(_3074_),
    .A3(_3078_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6474_ (.A1(_3003_),
    .A2(_2300_),
    .B1(_3004_),
    .B2(_2512_),
    .C1(_2518_),
    .C2(_3005_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6475_ (.A1(_3002_),
    .A2(_3080_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6476_ (.A1(_1676_),
    .A2(_3079_),
    .A3(_3081_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6477_ (.I(_2693_),
    .Z(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6478_ (.I(_2351_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6479_ (.A1(_2464_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][3] ),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6480_ (.A1(_3084_),
    .A2(_1855_),
    .B(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6481_ (.A1(_2635_),
    .A2(_3086_),
    .B(_1623_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6482_ (.A1(_2133_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][3] ),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6483_ (.A1(_2526_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][3] ),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6484_ (.A1(_2431_),
    .A2(_3088_),
    .A3(_3089_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6485_ (.A1(_3026_),
    .A2(_2502_),
    .B(_3090_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6486_ (.A1(_2066_),
    .A2(_2497_),
    .B(_3087_),
    .C(_3091_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6487_ (.A1(_3003_),
    .A2(_2306_),
    .B1(_3026_),
    .B2(_2485_),
    .C1(_2491_),
    .C2(_2499_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6488_ (.A1(_3002_),
    .A2(_3093_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6489_ (.A1(_3083_),
    .A2(_3092_),
    .A3(_3094_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6490_ (.A1(_3082_),
    .A2(_3095_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6491_ (.I(_2345_),
    .Z(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6492_ (.I0(\mod.Data_Mem.F_M.MRAM[12][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[14][4] ),
    .I2(\mod.Data_Mem.F_M.MRAM[13][4] ),
    .I3(_1870_),
    .S0(_2273_),
    .S1(_2500_),
    .Z(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6493_ (.A1(_2611_),
    .A2(\mod.Data_Mem.F_M.MRAM[1][4] ),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6494_ (.A1(_3084_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][4] ),
    .B(_2101_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6495_ (.A1(_2500_),
    .A2(\mod.Data_Mem.F_M.MRAM[2][4] ),
    .B(_2550_),
    .C(_2560_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6496_ (.A1(_3098_),
    .A2(_3099_),
    .B(_3100_),
    .ZN(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6497_ (.A1(_3096_),
    .A2(_3097_),
    .B(_3101_),
    .C(_2106_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6498_ (.A1(_3058_),
    .A2(_2549_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6499_ (.A1(_1623_),
    .A2(_3103_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6500_ (.A1(_3096_),
    .A2(_2313_),
    .B1(_2603_),
    .B2(_2546_),
    .C(_3104_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _6501_ (.I0(\mod.Data_Mem.F_M.MRAM[780][4] ),
    .I1(\mod.Data_Mem.F_M.MRAM[782][4] ),
    .I2(\mod.Data_Mem.F_M.MRAM[781][4] ),
    .I3(_1902_),
    .S0(_2264_),
    .S1(_2338_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6502_ (.A1(_3084_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][4] ),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6503_ (.A1(_2641_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][4] ),
    .B(_3058_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6504_ (.A1(_3107_),
    .A2(_3108_),
    .B(_2425_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6505_ (.A1(_2603_),
    .A2(_2537_),
    .B1(_3106_),
    .B2(_2204_),
    .C(_3109_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6506_ (.A1(_3047_),
    .A2(_2317_),
    .B1(_2488_),
    .B2(_2532_),
    .C1(_2530_),
    .C2(_2559_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6507_ (.A1(_3049_),
    .A2(_3111_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6508_ (.A1(_1491_),
    .A2(_3112_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6509_ (.A1(_3083_),
    .A2(_3102_),
    .A3(_3105_),
    .B1(_3110_),
    .B2(_3113_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6510_ (.A1(_2579_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][5] ),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6511_ (.I(_2374_),
    .Z(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6512_ (.A1(_2689_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][5] ),
    .B(_3115_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6513_ (.A1(_2075_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][5] ),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6514_ (.A1(_2418_),
    .A2(_1968_),
    .B(_2399_),
    .C(_3117_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6515_ (.A1(_3059_),
    .A2(_2583_),
    .B1(_2584_),
    .B2(_3019_),
    .C(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6516_ (.A1(_3114_),
    .A2(_3116_),
    .B(_3119_),
    .C(_3013_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6517_ (.A1(_3030_),
    .A2(_2323_),
    .B1(_3023_),
    .B2(_2569_),
    .C1(_2572_),
    .C2(_3022_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6518_ (.A1(_2827_),
    .A2(_3121_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6519_ (.A1(_3120_),
    .A2(_3122_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6520_ (.A1(_2641_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][5] ),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6521_ (.A1(_2558_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][5] ),
    .B(_3115_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6522_ (.A1(_2315_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][5] ),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6523_ (.A1(_2632_),
    .A2(_1955_),
    .B(_2399_),
    .C(_3126_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6524_ (.A1(_2488_),
    .A2(_2594_),
    .B(_3127_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6525_ (.A1(_2548_),
    .A2(_2589_),
    .B1(_3124_),
    .B2(_3125_),
    .C(_3128_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6526_ (.A1(_2203_),
    .A2(_2327_),
    .B1(_3059_),
    .B2(_2597_),
    .C1(_2598_),
    .C2(_3058_),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6527_ (.A1(_3049_),
    .A2(_3130_),
    .ZN(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6528_ (.A1(_2618_),
    .A2(_3129_),
    .B(_3131_),
    .C(_2073_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6529_ (.A1(_2523_),
    .A2(_3123_),
    .B(_3132_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6530_ (.A1(_2261_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][6] ),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6531_ (.A1(_2562_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][6] ),
    .B(_3115_),
    .C(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6532_ (.A1(_2289_),
    .A2(\mod.Data_Mem.F_M.MRAM[1][6] ),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6533_ (.A1(_2252_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][6] ),
    .B(_2100_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6534_ (.A1(_3135_),
    .A2(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6535_ (.A1(_3059_),
    .A2(_2636_),
    .B1(_2637_),
    .B2(_3019_),
    .C(_3137_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6536_ (.A1(_3013_),
    .A2(_3134_),
    .A3(_3138_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6537_ (.A1(_2065_),
    .A2(_2496_),
    .A3(_2628_),
    .B(_1758_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6538_ (.A1(_3096_),
    .A2(_2331_),
    .B1(_2623_),
    .B2(_3063_),
    .C(_3140_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6539_ (.A1(_2571_),
    .A2(\mod.Data_Mem.F_M.MRAM[781][6] ),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6540_ (.A1(_2611_),
    .A2(\mod.Data_Mem.F_M.MRAM[780][6] ),
    .B(_3142_),
    .C(_2168_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6541_ (.A1(_2089_),
    .A2(_2613_),
    .B(_3143_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6542_ (.A1(_3084_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][6] ),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6543_ (.A1(_2641_),
    .A2(\mod.Data_Mem.F_M.MRAM[769][6] ),
    .B(_2101_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6544_ (.A1(_3145_),
    .A2(_3146_),
    .B(_2425_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6545_ (.A1(_2603_),
    .A2(_2619_),
    .B1(_3144_),
    .B2(_2204_),
    .C(_3147_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6546_ (.A1(_3047_),
    .A2(_2334_),
    .B1(_2488_),
    .B2(_2607_),
    .C1(_2608_),
    .C2(_2559_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6547_ (.A1(_3049_),
    .A2(_3149_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6548_ (.A1(_1491_),
    .A2(_3150_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6549_ (.A1(_3083_),
    .A2(_3139_),
    .A3(_3141_),
    .B1(_3148_),
    .B2(_3151_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6550_ (.A1(_2722_),
    .A2(\mod.Data_Mem.F_M.MRAM[1][7] ),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6551_ (.A1(_2338_),
    .A2(\mod.Data_Mem.F_M.MRAM[0][7] ),
    .B(_2101_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6552_ (.A1(_2410_),
    .A2(\mod.Data_Mem.F_M.MRAM[12][7] ),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6553_ (.A1(_2722_),
    .A2(\mod.Data_Mem.F_M.MRAM[13][7] ),
    .B(_2387_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6554_ (.A1(_2538_),
    .A2(_2666_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6555_ (.A1(_3152_),
    .A2(_3153_),
    .B1(_3154_),
    .B2(_3155_),
    .C(_3156_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6556_ (.A1(_3020_),
    .A2(_2670_),
    .B(_3157_),
    .C(_2106_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6557_ (.A1(_2308_),
    .A2(_2496_),
    .A3(_2662_),
    .B(_1758_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6558_ (.A1(_3096_),
    .A2(_2340_),
    .B1(_2657_),
    .B2(_3063_),
    .C(_3159_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6559_ (.A1(_3030_),
    .A2(_2343_),
    .B1(_3023_),
    .B2(_2646_),
    .C1(_2644_),
    .C2(_2484_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6560_ (.A1(_2827_),
    .A2(_3161_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6561_ (.A1(\mod.Data_Mem.F_M.MRAM[781][7] ),
    .A2(_3115_),
    .B1(_3005_),
    .B2(\mod.Data_Mem.F_M.MRAM[769][7] ),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6562_ (.A1(_2391_),
    .A2(\mod.Data_Mem.F_M.MRAM[768][7] ),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6563_ (.A1(\mod.Data_Mem.F_M.MRAM[780][7] ),
    .A2(_1680_),
    .B1(_2559_),
    .B2(_3164_),
    .C(_2617_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6564_ (.A1(_2492_),
    .A2(_2649_),
    .B1(_2650_),
    .B2(_3008_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6565_ (.A1(_3016_),
    .A2(_3163_),
    .B(_3165_),
    .C(_3166_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6566_ (.A1(_2861_),
    .A2(_3162_),
    .A3(_3167_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6567_ (.A1(_3083_),
    .A2(_3158_),
    .A3(_3160_),
    .B(_3168_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6568_ (.I(\mod.I_addr[1] ),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6569_ (.A1(_0612_),
    .A2(_3169_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6570_ (.I(_3170_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6571_ (.I(\mod.I_addr[2] ),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6572_ (.A1(_0612_),
    .A2(_3169_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6573_ (.A1(_3171_),
    .A2(_3172_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6574_ (.I(_3173_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6575_ (.I(\mod.I_addr[3] ),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6576_ (.I(_3174_),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6577_ (.A1(\mod.I_addr[0] ),
    .A2(\mod.I_addr[2] ),
    .A3(\mod.I_addr[1] ),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6578_ (.A1(_3175_),
    .A2(_3176_),
    .Z(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6579_ (.I(_3177_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6580_ (.I(\mod.I_addr[4] ),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6581_ (.A1(_3175_),
    .A2(_3176_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6582_ (.A1(_3178_),
    .A2(_3179_),
    .Z(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6583_ (.I(_3180_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6584_ (.A1(_3178_),
    .A2(_3179_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6585_ (.A1(\mod.I_addr[5] ),
    .A2(_3181_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6586_ (.I(_3182_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6587_ (.A1(_3178_),
    .A2(\mod.I_addr[5] ),
    .A3(_3179_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6588_ (.A1(\mod.I_addr[6] ),
    .A2(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6589_ (.I(_3184_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6590_ (.A1(_3178_),
    .A2(\mod.I_addr[6] ),
    .A3(\mod.I_addr[5] ),
    .A4(_3179_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6591_ (.A1(\mod.I_addr[7] ),
    .A2(_3185_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6592_ (.I(_3186_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6593_ (.I(\mod.Data_Mem.F_M.MRAM[11][0] ),
    .Z(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6594_ (.I(_3187_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6595_ (.I(\mod.Data_Mem.F_M.MRAM[11][1] ),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6596_ (.I(_3188_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6597_ (.I(\mod.Data_Mem.F_M.MRAM[11][2] ),
    .Z(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6598_ (.I(_3189_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6599_ (.I(\mod.Data_Mem.F_M.MRAM[11][3] ),
    .Z(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6600_ (.I(_3190_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6601_ (.I(\mod.Data_Mem.F_M.MRAM[11][4] ),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6602_ (.I(_3191_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6603_ (.I(\mod.Data_Mem.F_M.MRAM[11][5] ),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6604_ (.I(_3192_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6605_ (.I(\mod.Data_Mem.F_M.MRAM[11][6] ),
    .Z(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6606_ (.I(_3193_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6607_ (.I(\mod.Data_Mem.F_M.MRAM[11][7] ),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6608_ (.I(_3194_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6609_ (.I(\mod.Data_Mem.F_M.MRAM[24][0] ),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6610_ (.I(_3195_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6611_ (.I(\mod.Data_Mem.F_M.MRAM[24][1] ),
    .Z(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6612_ (.I(_3196_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6613_ (.I(\mod.Data_Mem.F_M.MRAM[24][2] ),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6614_ (.I(_3197_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6615_ (.I(\mod.Data_Mem.F_M.MRAM[24][3] ),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6616_ (.I(_3198_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6617_ (.I(\mod.Data_Mem.F_M.MRAM[24][4] ),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6618_ (.I(_3199_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6619_ (.I(\mod.Data_Mem.F_M.MRAM[24][5] ),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6620_ (.I(_3200_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6621_ (.I(\mod.Data_Mem.F_M.MRAM[24][6] ),
    .Z(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6622_ (.I(_3201_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6623_ (.I(\mod.Data_Mem.F_M.MRAM[24][7] ),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6624_ (.I(_3202_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6625_ (.I(\mod.Data_Mem.F_M.MRAM[26][0] ),
    .Z(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6626_ (.I(_3203_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6627_ (.I(\mod.Data_Mem.F_M.MRAM[26][1] ),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6628_ (.I(_3204_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6629_ (.I(\mod.Data_Mem.F_M.MRAM[26][2] ),
    .Z(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6630_ (.I(_3205_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6631_ (.I(\mod.Data_Mem.F_M.MRAM[26][3] ),
    .Z(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6632_ (.I(_3206_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6633_ (.I(\mod.Data_Mem.F_M.MRAM[26][4] ),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6634_ (.I(_3207_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6635_ (.I(\mod.Data_Mem.F_M.MRAM[26][5] ),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6636_ (.I(_3208_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6637_ (.I(\mod.Data_Mem.F_M.MRAM[26][6] ),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6638_ (.I(_3209_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6639_ (.I(\mod.Data_Mem.F_M.MRAM[26][7] ),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6640_ (.I(_3210_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6641_ (.I(\mod.Data_Mem.F_M.MRAM[25][0] ),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6642_ (.I(_3211_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6643_ (.I(\mod.Data_Mem.F_M.MRAM[25][1] ),
    .Z(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6644_ (.I(_3212_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6645_ (.I(\mod.Data_Mem.F_M.MRAM[25][2] ),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6646_ (.I(_3213_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6647_ (.I(\mod.Data_Mem.F_M.MRAM[25][3] ),
    .Z(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6648_ (.I(_3214_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6649_ (.I(\mod.Data_Mem.F_M.MRAM[25][4] ),
    .Z(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6650_ (.I(_3215_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6651_ (.I(\mod.Data_Mem.F_M.MRAM[25][5] ),
    .Z(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6652_ (.I(_3216_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6653_ (.I(\mod.Data_Mem.F_M.MRAM[25][6] ),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6654_ (.I(_3217_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6655_ (.I(\mod.Data_Mem.F_M.MRAM[25][7] ),
    .Z(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6656_ (.I(_3218_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6657_ (.I(\mod.Data_Mem.F_M.MRAM[27][0] ),
    .Z(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6658_ (.I(_3219_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6659_ (.I(\mod.Data_Mem.F_M.MRAM[27][1] ),
    .Z(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6660_ (.I(_3220_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6661_ (.I(\mod.Data_Mem.F_M.MRAM[27][2] ),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6662_ (.I(_3221_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6663_ (.I(\mod.Data_Mem.F_M.MRAM[27][3] ),
    .Z(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6664_ (.I(_3222_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6665_ (.I(\mod.Data_Mem.F_M.MRAM[27][4] ),
    .Z(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6666_ (.I(_3223_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6667_ (.I(\mod.Data_Mem.F_M.MRAM[27][5] ),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6668_ (.I(_3224_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6669_ (.I(\mod.Data_Mem.F_M.MRAM[27][6] ),
    .Z(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6670_ (.I(_3225_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6671_ (.I(\mod.Data_Mem.F_M.MRAM[27][7] ),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6672_ (.I(_3226_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6673_ (.I(net3),
    .Z(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6674_ (.I(_3227_),
    .Z(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6675_ (.A1(\mod.Data_Mem.F_M.dest[4] ),
    .A2(\mod.Data_Mem.F_M.dest[2] ),
    .Z(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6676_ (.I(_3229_),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6677_ (.A1(\mod.Data_Mem.F_M.dest[1] ),
    .A2(\mod.Data_Mem.F_M.dest[0] ),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6678_ (.I(_3231_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6679_ (.I(\mod.DMen_reg2 ),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6680_ (.A1(\mod.Data_Mem.F_M.dest[8] ),
    .A2(_3233_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6681_ (.I(_3234_),
    .Z(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6682_ (.A1(_3230_),
    .A2(_3232_),
    .A3(_3235_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6683_ (.I(_3236_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6684_ (.I0(_3228_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][0] ),
    .S(_3237_),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6685_ (.I(_3238_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6686_ (.I(net4),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6687_ (.I(_3239_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6688_ (.I0(_3240_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][1] ),
    .S(_3237_),
    .Z(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6689_ (.I(_3241_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6690_ (.I(net5),
    .Z(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6691_ (.I(_3242_),
    .Z(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6692_ (.I0(_3243_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][2] ),
    .S(_3237_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6693_ (.I(_3244_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6694_ (.I(net6),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6695_ (.I(_3245_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6696_ (.I0(_3246_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][3] ),
    .S(_3237_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6697_ (.I(_3247_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6698_ (.I(net7),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6699_ (.I(_3248_),
    .Z(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6700_ (.I(_3236_),
    .Z(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6701_ (.I0(_3249_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][4] ),
    .S(_3250_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6702_ (.I(_3251_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6703_ (.I(net8),
    .Z(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6704_ (.I(_3252_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6705_ (.I0(_3253_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][5] ),
    .S(_3250_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6706_ (.I(_3254_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6707_ (.I(net9),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6708_ (.I(_3255_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6709_ (.I0(_3256_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][6] ),
    .S(_3250_),
    .Z(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6710_ (.I(_3257_),
    .Z(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6711_ (.I(net10),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6712_ (.I(_3258_),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6713_ (.I0(_3259_),
    .I1(\mod.Data_Mem.F_M.MRAM[28][7] ),
    .S(_3250_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6714_ (.I(_3260_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6715_ (.I(\mod.Data_Mem.F_M.MRAM[10][0] ),
    .Z(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6716_ (.I(_3261_),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6717_ (.I(\mod.Data_Mem.F_M.MRAM[10][1] ),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6718_ (.I(_3262_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6719_ (.I(\mod.Data_Mem.F_M.MRAM[10][2] ),
    .Z(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6720_ (.I(_3263_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6721_ (.I(\mod.Data_Mem.F_M.MRAM[10][3] ),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6722_ (.I(_3264_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6723_ (.I(\mod.Data_Mem.F_M.MRAM[10][4] ),
    .Z(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6724_ (.I(_3265_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6725_ (.I(\mod.Data_Mem.F_M.MRAM[10][5] ),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6726_ (.I(_3266_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6727_ (.I(\mod.Data_Mem.F_M.MRAM[10][6] ),
    .Z(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6728_ (.I(_3267_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6729_ (.I(\mod.Data_Mem.F_M.MRAM[10][7] ),
    .Z(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6730_ (.I(_3268_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6731_ (.I(_3231_),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6732_ (.I(_3234_),
    .Z(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6733_ (.A1(\mod.Data_Mem.F_M.dest[4] ),
    .A2(\mod.Data_Mem.F_M.dest[2] ),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6734_ (.I(_3271_),
    .Z(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6735_ (.A1(_3269_),
    .A2(_3270_),
    .A3(_3272_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6736_ (.I(_3273_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6737_ (.I0(_3228_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][0] ),
    .S(_3274_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6738_ (.I(_3275_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6739_ (.I0(_3240_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][1] ),
    .S(_3274_),
    .Z(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6740_ (.I(_3276_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6741_ (.I0(_3243_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][2] ),
    .S(_3274_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6742_ (.I(_3277_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6743_ (.I0(_3246_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][3] ),
    .S(_3274_),
    .Z(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6744_ (.I(_3278_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6745_ (.I(_3273_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6746_ (.I0(_3249_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][4] ),
    .S(_3279_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6747_ (.I(_3280_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6748_ (.I0(_3253_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][5] ),
    .S(_3279_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6749_ (.I(_3281_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6750_ (.I0(_3256_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][6] ),
    .S(_3279_),
    .Z(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6751_ (.I(_3282_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6752_ (.I0(_3259_),
    .I1(\mod.Data_Mem.F_M.MRAM[0][7] ),
    .S(_3279_),
    .Z(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6753_ (.I(_3283_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6754_ (.I(\mod.Data_Mem.F_M.MRAM[8][0] ),
    .Z(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6755_ (.I(_3284_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6756_ (.I(\mod.Data_Mem.F_M.MRAM[8][1] ),
    .Z(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6757_ (.I(_3285_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6758_ (.I(\mod.Data_Mem.F_M.MRAM[8][2] ),
    .Z(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6759_ (.I(_3286_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6760_ (.I(\mod.Data_Mem.F_M.MRAM[8][3] ),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6761_ (.I(_3287_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6762_ (.I(\mod.Data_Mem.F_M.MRAM[8][4] ),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6763_ (.I(_3288_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6764_ (.I(\mod.Data_Mem.F_M.MRAM[8][5] ),
    .Z(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6765_ (.I(_3289_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6766_ (.I(\mod.Data_Mem.F_M.MRAM[8][6] ),
    .Z(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6767_ (.I(_3290_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6768_ (.I(\mod.Data_Mem.F_M.MRAM[8][7] ),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6769_ (.I(_3291_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6770_ (.I(net3),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6771_ (.I(_3292_),
    .Z(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6772_ (.I(_3229_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6773_ (.A1(\mod.Data_Mem.F_M.dest[1] ),
    .A2(\mod.Data_Mem.F_M.dest[0] ),
    .Z(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6774_ (.I(_3295_),
    .Z(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6775_ (.A1(\mod.Data_Mem.F_M.dest[8] ),
    .A2(\mod.DMen_reg2 ),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6776_ (.I(_3297_),
    .Z(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6777_ (.A1(_3294_),
    .A2(_3296_),
    .A3(_3298_),
    .Z(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6778_ (.I(_3299_),
    .Z(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6779_ (.I0(\mod.Data_Mem.F_M.MRAM[799][0] ),
    .I1(_3293_),
    .S(_3300_),
    .Z(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6780_ (.I(_3301_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6781_ (.I(net4),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6782_ (.I(_3302_),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6783_ (.I0(\mod.Data_Mem.F_M.MRAM[799][1] ),
    .I1(_3303_),
    .S(_3300_),
    .Z(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6784_ (.I(_3304_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6785_ (.I(net5),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6786_ (.I(_3305_),
    .Z(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6787_ (.I0(\mod.Data_Mem.F_M.MRAM[799][2] ),
    .I1(_3306_),
    .S(_3300_),
    .Z(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6788_ (.I(_3307_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6789_ (.I(net6),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6790_ (.I(_3308_),
    .Z(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6791_ (.I0(\mod.Data_Mem.F_M.MRAM[799][3] ),
    .I1(_3309_),
    .S(_3300_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6792_ (.I(_3310_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6793_ (.I(net7),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6794_ (.I(_3311_),
    .Z(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6795_ (.I(_3299_),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6796_ (.I0(\mod.Data_Mem.F_M.MRAM[799][4] ),
    .I1(_3312_),
    .S(_3313_),
    .Z(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6797_ (.I(_3314_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6798_ (.I(net8),
    .Z(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6799_ (.I(_3315_),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6800_ (.I0(\mod.Data_Mem.F_M.MRAM[799][5] ),
    .I1(_3316_),
    .S(_3313_),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6801_ (.I(_3317_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6802_ (.I(net9),
    .Z(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6803_ (.I(_3318_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6804_ (.I0(\mod.Data_Mem.F_M.MRAM[799][6] ),
    .I1(_3319_),
    .S(_3313_),
    .Z(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6805_ (.I(_3320_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6806_ (.I(net10),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6807_ (.I(_3321_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6808_ (.I0(\mod.Data_Mem.F_M.MRAM[799][7] ),
    .I1(_3322_),
    .S(_3313_),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6809_ (.I(_3323_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6810_ (.I(\mod.Data_Mem.F_M.MRAM[789][0] ),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6811_ (.I(_3324_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6812_ (.I(\mod.Data_Mem.F_M.MRAM[789][1] ),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6813_ (.I(_3325_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6814_ (.I(\mod.Data_Mem.F_M.MRAM[789][2] ),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6815_ (.I(_3326_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6816_ (.I(\mod.Data_Mem.F_M.MRAM[789][3] ),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6817_ (.I(_3327_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6818_ (.I(\mod.Data_Mem.F_M.MRAM[789][4] ),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6819_ (.I(_3328_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6820_ (.I(\mod.Data_Mem.F_M.MRAM[789][5] ),
    .Z(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6821_ (.I(_3329_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6822_ (.I(\mod.Data_Mem.F_M.MRAM[789][6] ),
    .Z(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6823_ (.I(_3330_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6824_ (.I(\mod.Data_Mem.F_M.MRAM[789][7] ),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6825_ (.I(_3331_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6826_ (.I(_3271_),
    .Z(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6827_ (.I(\mod.Data_Mem.F_M.dest[0] ),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6828_ (.A1(\mod.Data_Mem.F_M.dest[1] ),
    .A2(_3333_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6829_ (.I(_3334_),
    .Z(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6830_ (.A1(_3332_),
    .A2(_3298_),
    .A3(_3335_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6831_ (.I(_3336_),
    .Z(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6832_ (.I0(_3228_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][0] ),
    .S(_3337_),
    .Z(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6833_ (.I(_3338_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6834_ (.I0(_3240_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][1] ),
    .S(_3337_),
    .Z(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6835_ (.I(_3339_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6836_ (.I(_3336_),
    .Z(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6837_ (.I0(_3243_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][2] ),
    .S(_3340_),
    .Z(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6838_ (.I(_3341_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6839_ (.I0(_3246_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][3] ),
    .S(_3340_),
    .Z(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6840_ (.I(_3342_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6841_ (.I0(_3249_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][4] ),
    .S(_3340_),
    .Z(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6842_ (.I(_3343_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6843_ (.A1(_3316_),
    .A2(_3337_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6844_ (.A1(_1955_),
    .A2(_3337_),
    .B(_3344_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6845_ (.I0(_3256_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][6] ),
    .S(_3340_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6846_ (.I(_3345_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6847_ (.I0(_3259_),
    .I1(\mod.Data_Mem.F_M.MRAM[769][7] ),
    .S(_3336_),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6848_ (.I(_3346_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6849_ (.I(\mod.Data_Mem.F_M.MRAM[779][0] ),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6850_ (.I(_3347_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6851_ (.I(\mod.Data_Mem.F_M.MRAM[779][1] ),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6852_ (.I(_3348_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6853_ (.I(\mod.Data_Mem.F_M.MRAM[779][2] ),
    .Z(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6854_ (.I(_3349_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6855_ (.I(\mod.Data_Mem.F_M.MRAM[779][3] ),
    .Z(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6856_ (.I(_3350_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6857_ (.I(\mod.Data_Mem.F_M.MRAM[779][4] ),
    .Z(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6858_ (.I(_3351_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6859_ (.I(\mod.Data_Mem.F_M.MRAM[779][5] ),
    .Z(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6860_ (.I(_3352_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6861_ (.I(\mod.Data_Mem.F_M.MRAM[779][6] ),
    .Z(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6862_ (.I(_3353_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6863_ (.I(\mod.Data_Mem.F_M.MRAM[779][7] ),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6864_ (.I(_3354_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6865_ (.I(\mod.Data_Mem.F_M.MRAM[6][0] ),
    .Z(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6866_ (.I(_3355_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6867_ (.I(\mod.Data_Mem.F_M.MRAM[6][1] ),
    .Z(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6868_ (.I(_3356_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6869_ (.I(\mod.Data_Mem.F_M.MRAM[6][2] ),
    .Z(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6870_ (.I(_3357_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6871_ (.I(\mod.Data_Mem.F_M.MRAM[6][3] ),
    .Z(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6872_ (.I(_3358_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6873_ (.I(\mod.Data_Mem.F_M.MRAM[6][4] ),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6874_ (.I(_3359_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6875_ (.I(\mod.Data_Mem.F_M.MRAM[6][5] ),
    .Z(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6876_ (.I(_3360_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6877_ (.I(\mod.Data_Mem.F_M.MRAM[6][6] ),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6878_ (.I(_3361_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6879_ (.I(\mod.Data_Mem.F_M.MRAM[6][7] ),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6880_ (.I(_3362_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6881_ (.I(\mod.Data_Mem.F_M.MRAM[4][0] ),
    .Z(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6882_ (.I(_3363_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6883_ (.I(\mod.Data_Mem.F_M.MRAM[4][1] ),
    .Z(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6884_ (.I(_3364_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6885_ (.I(\mod.Data_Mem.F_M.MRAM[4][2] ),
    .Z(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6886_ (.I(_3365_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6887_ (.I(\mod.Data_Mem.F_M.MRAM[4][3] ),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6888_ (.I(_3366_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6889_ (.I(\mod.Data_Mem.F_M.MRAM[4][4] ),
    .Z(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6890_ (.I(_3367_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6891_ (.I(\mod.Data_Mem.F_M.MRAM[4][5] ),
    .Z(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6892_ (.I(_3368_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6893_ (.I(\mod.Data_Mem.F_M.MRAM[4][6] ),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6894_ (.I(_3369_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6895_ (.I(\mod.Data_Mem.F_M.MRAM[4][7] ),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6896_ (.I(_3370_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6897_ (.I(_3334_),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6898_ (.I(\mod.Data_Mem.F_M.dest[2] ),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6899_ (.A1(\mod.Data_Mem.F_M.dest[4] ),
    .A2(_3372_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6900_ (.I(_3373_),
    .Z(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6901_ (.A1(_3235_),
    .A2(_3371_),
    .A3(_3374_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6902_ (.I(_3375_),
    .Z(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6903_ (.I0(_3228_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][0] ),
    .S(_3376_),
    .Z(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6904_ (.I(_3377_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6905_ (.I0(_3240_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][1] ),
    .S(_3376_),
    .Z(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6906_ (.I(_3378_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6907_ (.I0(_3243_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][2] ),
    .S(_3376_),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6908_ (.I(_3379_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6909_ (.I0(_3246_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][3] ),
    .S(_3376_),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6910_ (.I(_3380_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6911_ (.I(_3375_),
    .Z(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6912_ (.I0(_3249_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][4] ),
    .S(_3381_),
    .Z(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6913_ (.I(_3382_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6914_ (.I0(_3253_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][5] ),
    .S(_3381_),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6915_ (.I(_3383_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6916_ (.I0(_3256_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][6] ),
    .S(_3381_),
    .Z(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6917_ (.I(_3384_),
    .Z(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6918_ (.I0(_3259_),
    .I1(\mod.Data_Mem.F_M.MRAM[13][7] ),
    .S(_3381_),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6919_ (.I(_3385_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6920_ (.I(_3227_),
    .Z(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6921_ (.I(_3373_),
    .Z(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6922_ (.A1(\mod.Data_Mem.F_M.dest[1] ),
    .A2(_3333_),
    .Z(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6923_ (.I(_3388_),
    .Z(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6924_ (.A1(_3235_),
    .A2(_3387_),
    .A3(_3389_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6925_ (.I(_3390_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6926_ (.I0(_3386_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][0] ),
    .S(_3391_),
    .Z(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6927_ (.I(_3392_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6928_ (.I(_3239_),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6929_ (.I0(_3393_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][1] ),
    .S(_3391_),
    .Z(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6930_ (.I(_3394_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6931_ (.I(_3242_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6932_ (.I0(_3395_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][2] ),
    .S(_3391_),
    .Z(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6933_ (.I(_3396_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6934_ (.I(_3245_),
    .Z(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6935_ (.I0(_3397_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][3] ),
    .S(_3391_),
    .Z(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6936_ (.I(_3398_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6937_ (.I(_3248_),
    .Z(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6938_ (.I(_3390_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6939_ (.I0(_3399_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][4] ),
    .S(_3400_),
    .Z(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6940_ (.I(_3401_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6941_ (.I0(_3253_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][5] ),
    .S(_3400_),
    .Z(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6942_ (.I(_3402_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6943_ (.I(_3255_),
    .Z(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6944_ (.I0(_3403_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][6] ),
    .S(_3400_),
    .Z(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6945_ (.I(_3404_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6946_ (.I(_3258_),
    .Z(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6947_ (.I0(_3405_),
    .I1(\mod.Data_Mem.F_M.MRAM[14][7] ),
    .S(_3400_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6948_ (.I(_3406_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6949_ (.I(_3295_),
    .Z(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6950_ (.A1(_3235_),
    .A2(_3407_),
    .A3(_3374_),
    .ZN(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6951_ (.I(_3408_),
    .Z(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6952_ (.I0(_3386_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][0] ),
    .S(_3409_),
    .Z(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6953_ (.I(_3410_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6954_ (.I0(_3393_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][1] ),
    .S(_3409_),
    .Z(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6955_ (.I(_3411_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6956_ (.I0(_3395_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][2] ),
    .S(_3409_),
    .Z(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6957_ (.I(_3412_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6958_ (.I0(_3397_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][3] ),
    .S(_3409_),
    .Z(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6959_ (.I(_3413_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6960_ (.I(_3408_),
    .Z(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6961_ (.I0(_3399_),
    .I1(_1870_),
    .S(_3414_),
    .Z(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6962_ (.I(_3415_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6963_ (.I(_3252_),
    .Z(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6964_ (.I0(_3416_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][5] ),
    .S(_3414_),
    .Z(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6965_ (.I(_3417_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6966_ (.I0(_3403_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][6] ),
    .S(_3414_),
    .Z(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6967_ (.I(_3418_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6968_ (.I0(_3405_),
    .I1(\mod.Data_Mem.F_M.MRAM[15][7] ),
    .S(_3414_),
    .Z(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6969_ (.I(_3419_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6970_ (.A1(\mod.Data_Mem.F_M.dest[4] ),
    .A2(_3372_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6971_ (.I(_3420_),
    .Z(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6972_ (.A1(_3269_),
    .A2(_3270_),
    .A3(_3421_),
    .ZN(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6973_ (.I(_3422_),
    .Z(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6974_ (.I0(_3386_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][0] ),
    .S(_3423_),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6975_ (.I(_3424_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6976_ (.I0(_3393_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][1] ),
    .S(_3423_),
    .Z(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6977_ (.I(_3425_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6978_ (.I0(_3395_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][2] ),
    .S(_3423_),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6979_ (.I(_3426_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6980_ (.I0(_3397_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][3] ),
    .S(_3423_),
    .Z(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6981_ (.I(_3427_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6982_ (.I(_3422_),
    .Z(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6983_ (.I0(_3399_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][4] ),
    .S(_3428_),
    .Z(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6984_ (.I(_3429_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6985_ (.I0(_3416_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][5] ),
    .S(_3428_),
    .Z(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6986_ (.I(_3430_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6987_ (.I0(_3403_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][6] ),
    .S(_3428_),
    .Z(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6988_ (.I(_3431_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6989_ (.I0(_3405_),
    .I1(\mod.Data_Mem.F_M.MRAM[16][7] ),
    .S(_3428_),
    .Z(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6990_ (.I(_3432_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6991_ (.I(_3234_),
    .Z(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6992_ (.A1(_3433_),
    .A2(_3371_),
    .A3(_3421_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6993_ (.I(_3434_),
    .Z(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6994_ (.I0(_3386_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][0] ),
    .S(_3435_),
    .Z(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6995_ (.I(_3436_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6996_ (.I0(_3393_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][1] ),
    .S(_3435_),
    .Z(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6997_ (.I(_3437_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6998_ (.I0(_3395_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][2] ),
    .S(_3435_),
    .Z(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6999_ (.I(_3438_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7000_ (.I0(_3397_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][3] ),
    .S(_3435_),
    .Z(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7001_ (.I(_3439_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7002_ (.I(_3434_),
    .Z(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7003_ (.I0(_3399_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][4] ),
    .S(_3440_),
    .Z(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7004_ (.I(_3441_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7005_ (.I0(_3416_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][5] ),
    .S(_3440_),
    .Z(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7006_ (.I(_3442_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7007_ (.I0(_3403_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][6] ),
    .S(_3440_),
    .Z(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7008_ (.I(_3443_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7009_ (.I0(_3405_),
    .I1(\mod.Data_Mem.F_M.MRAM[17][7] ),
    .S(_3440_),
    .Z(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7010_ (.I(_3444_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7011_ (.I(_3227_),
    .Z(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7012_ (.I(_3388_),
    .Z(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7013_ (.A1(_3433_),
    .A2(_3446_),
    .A3(_3421_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7014_ (.I(_3447_),
    .Z(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7015_ (.I0(_3445_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][0] ),
    .S(_3448_),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7016_ (.I(_3449_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7017_ (.I(_3239_),
    .Z(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7018_ (.I0(_3450_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][1] ),
    .S(_3448_),
    .Z(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7019_ (.I(_3451_),
    .Z(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7020_ (.I(_3242_),
    .Z(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7021_ (.I0(_3452_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][2] ),
    .S(_3448_),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7022_ (.I(_3453_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7023_ (.I(_3245_),
    .Z(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7024_ (.I0(_3454_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][3] ),
    .S(_3448_),
    .Z(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7025_ (.I(_3455_),
    .Z(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7026_ (.I(_3248_),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7027_ (.I(_3447_),
    .Z(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7028_ (.I0(_3456_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][4] ),
    .S(_3457_),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7029_ (.I(_3458_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7030_ (.I0(_3416_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][5] ),
    .S(_3457_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7031_ (.I(_3459_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7032_ (.I(_3255_),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7033_ (.I0(_3460_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][6] ),
    .S(_3457_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7034_ (.I(_3461_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7035_ (.I(_3258_),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7036_ (.I0(_3462_),
    .I1(\mod.Data_Mem.F_M.MRAM[18][7] ),
    .S(_3457_),
    .Z(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7037_ (.I(_3463_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7038_ (.I(_3234_),
    .Z(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7039_ (.A1(_3464_),
    .A2(_3332_),
    .A3(_3335_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7040_ (.I(_3465_),
    .Z(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7041_ (.I0(_3445_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][0] ),
    .S(_3466_),
    .Z(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7042_ (.I(_3467_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7043_ (.I0(_3450_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][1] ),
    .S(_3466_),
    .Z(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7044_ (.I(_3468_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7045_ (.I(_3465_),
    .Z(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7046_ (.I0(_3452_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][2] ),
    .S(_3469_),
    .Z(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7047_ (.I(_3470_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7048_ (.I0(_3454_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][3] ),
    .S(_3469_),
    .Z(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7049_ (.I(_3471_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7050_ (.I0(_3456_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][4] ),
    .S(_3469_),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7051_ (.I(_3472_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7052_ (.A1(_3316_),
    .A2(_3466_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7053_ (.A1(_1968_),
    .A2(_3466_),
    .B(_3473_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7054_ (.I0(_3460_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][6] ),
    .S(_3469_),
    .Z(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7055_ (.I(_3474_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7056_ (.I0(_3462_),
    .I1(\mod.Data_Mem.F_M.MRAM[1][7] ),
    .S(_3465_),
    .Z(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7057_ (.I(_3475_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7058_ (.I(\mod.Data_Mem.F_M.MRAM[20][0] ),
    .Z(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7059_ (.I(_3476_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7060_ (.I(\mod.Data_Mem.F_M.MRAM[20][1] ),
    .Z(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7061_ (.I(_3477_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7062_ (.I(\mod.Data_Mem.F_M.MRAM[20][2] ),
    .Z(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7063_ (.I(_3478_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7064_ (.I(\mod.Data_Mem.F_M.MRAM[20][3] ),
    .Z(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7065_ (.I(_3479_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7066_ (.I(\mod.Data_Mem.F_M.MRAM[20][4] ),
    .Z(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7067_ (.I(_3480_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7068_ (.I(\mod.Data_Mem.F_M.MRAM[20][5] ),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7069_ (.I(_3481_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7070_ (.I(\mod.Data_Mem.F_M.MRAM[20][6] ),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7071_ (.I(_3482_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7072_ (.I(\mod.Data_Mem.F_M.MRAM[20][7] ),
    .Z(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7073_ (.I(_3483_),
    .Z(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7074_ (.I(\mod.Data_Mem.F_M.MRAM[21][0] ),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7075_ (.I(_3484_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7076_ (.I(\mod.Data_Mem.F_M.MRAM[21][1] ),
    .Z(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7077_ (.I(_3485_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7078_ (.I(\mod.Data_Mem.F_M.MRAM[21][2] ),
    .Z(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7079_ (.I(_3486_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7080_ (.I(\mod.Data_Mem.F_M.MRAM[21][3] ),
    .Z(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7081_ (.I(_3487_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7082_ (.I(\mod.Data_Mem.F_M.MRAM[21][4] ),
    .Z(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7083_ (.I(_3488_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7084_ (.I(\mod.Data_Mem.F_M.MRAM[21][5] ),
    .Z(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7085_ (.I(_3489_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7086_ (.I(\mod.Data_Mem.F_M.MRAM[21][6] ),
    .Z(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7087_ (.I(_3490_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7088_ (.I(\mod.Data_Mem.F_M.MRAM[21][7] ),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7089_ (.I(_3491_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7090_ (.I(\mod.Data_Mem.F_M.MRAM[23][0] ),
    .Z(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7091_ (.I(_3492_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7092_ (.I(\mod.Data_Mem.F_M.MRAM[23][1] ),
    .Z(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7093_ (.I(_3493_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7094_ (.I(\mod.Data_Mem.F_M.MRAM[23][2] ),
    .Z(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7095_ (.I(_3494_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7096_ (.I(\mod.Data_Mem.F_M.MRAM[23][3] ),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7097_ (.I(_3495_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7098_ (.I(\mod.Data_Mem.F_M.MRAM[23][4] ),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7099_ (.I(_3496_),
    .Z(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7100_ (.I(\mod.Data_Mem.F_M.MRAM[23][5] ),
    .Z(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7101_ (.I(_3497_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7102_ (.I(\mod.Data_Mem.F_M.MRAM[23][6] ),
    .Z(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7103_ (.I(_3498_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7104_ (.I(\mod.Data_Mem.F_M.MRAM[23][7] ),
    .Z(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7105_ (.I(_3499_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7106_ (.A1(_3433_),
    .A2(_3272_),
    .A3(_3407_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7107_ (.I(_3500_),
    .Z(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7108_ (.I0(_3445_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][0] ),
    .S(_3501_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7109_ (.I(_3502_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7110_ (.I0(_3450_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][1] ),
    .S(_3501_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7111_ (.I(_3503_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7112_ (.I0(_3452_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][2] ),
    .S(_3501_),
    .Z(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7113_ (.I(_3504_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7114_ (.I0(_3454_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][3] ),
    .S(_3501_),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7115_ (.I(_3505_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7116_ (.I(_3500_),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7117_ (.I0(_3456_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][4] ),
    .S(_3506_),
    .Z(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7118_ (.I(_3507_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7119_ (.I(_3252_),
    .Z(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7120_ (.I0(_3508_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][5] ),
    .S(_3506_),
    .Z(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7121_ (.I(_3509_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7122_ (.I0(_3460_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][6] ),
    .S(_3506_),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7123_ (.I(_3510_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7124_ (.I0(_3462_),
    .I1(\mod.Data_Mem.F_M.MRAM[3][7] ),
    .S(_3506_),
    .Z(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7125_ (.I(_3511_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7126_ (.A1(_3433_),
    .A2(_3407_),
    .A3(_3421_),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7127_ (.I(_3512_),
    .Z(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7128_ (.I0(_3445_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][0] ),
    .S(_3513_),
    .Z(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7129_ (.I(_3514_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7130_ (.I0(_3450_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][1] ),
    .S(_3513_),
    .Z(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7131_ (.I(_3515_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7132_ (.I0(_3452_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][2] ),
    .S(_3513_),
    .Z(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7133_ (.I(_3516_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7134_ (.I0(_3454_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][3] ),
    .S(_3513_),
    .Z(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7135_ (.I(_3517_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7136_ (.I(_3512_),
    .Z(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7137_ (.I0(_3456_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][4] ),
    .S(_3518_),
    .Z(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7138_ (.I(_3519_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7139_ (.I0(_3508_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][5] ),
    .S(_3518_),
    .Z(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7140_ (.I(_3520_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7141_ (.I0(_3460_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][6] ),
    .S(_3518_),
    .Z(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7142_ (.I(_3521_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7143_ (.I0(_3462_),
    .I1(\mod.Data_Mem.F_M.MRAM[19][7] ),
    .S(_3518_),
    .Z(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7144_ (.I(_3522_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7145_ (.I(_3227_),
    .Z(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7146_ (.A1(_3269_),
    .A2(_3270_),
    .A3(_3374_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7147_ (.I(_3524_),
    .Z(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7148_ (.I0(_3523_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][0] ),
    .S(_3525_),
    .Z(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7149_ (.I(_3526_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7150_ (.I(_3239_),
    .Z(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7151_ (.I0(_3527_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][1] ),
    .S(_3525_),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7152_ (.I(_3528_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7153_ (.I(_3242_),
    .Z(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7154_ (.I0(_3529_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][2] ),
    .S(_3525_),
    .Z(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7155_ (.I(_3530_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7156_ (.I(_3245_),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7157_ (.I0(_3531_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][3] ),
    .S(_3525_),
    .Z(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7158_ (.I(_3532_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7159_ (.I(_3248_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7160_ (.I(_3524_),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7161_ (.I0(_3533_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][4] ),
    .S(_3534_),
    .Z(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7162_ (.I(_3535_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7163_ (.I0(_3508_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][5] ),
    .S(_3534_),
    .Z(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7164_ (.I(_3536_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7165_ (.I(_3255_),
    .Z(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7166_ (.I0(_3537_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][6] ),
    .S(_3534_),
    .Z(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7167_ (.I(_3538_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7168_ (.I(_3258_),
    .Z(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7169_ (.I0(_3539_),
    .I1(\mod.Data_Mem.F_M.MRAM[12][7] ),
    .S(_3534_),
    .Z(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7170_ (.I(_3540_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7171_ (.I(\mod.Data_Mem.F_M.MRAM[22][0] ),
    .Z(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7172_ (.I(_3541_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7173_ (.I(\mod.Data_Mem.F_M.MRAM[22][1] ),
    .Z(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7174_ (.I(_3542_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7175_ (.I(\mod.Data_Mem.F_M.MRAM[22][2] ),
    .Z(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7176_ (.I(_3543_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7177_ (.I(\mod.Data_Mem.F_M.MRAM[22][3] ),
    .Z(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7178_ (.I(_3544_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7179_ (.I(\mod.Data_Mem.F_M.MRAM[22][4] ),
    .Z(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7180_ (.I(_3545_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7181_ (.I(\mod.Data_Mem.F_M.MRAM[22][5] ),
    .Z(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7182_ (.I(_3546_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7183_ (.I(\mod.Data_Mem.F_M.MRAM[22][6] ),
    .Z(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7184_ (.I(_3547_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7185_ (.I(\mod.Data_Mem.F_M.MRAM[22][7] ),
    .Z(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7186_ (.I(_3548_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7187_ (.A1(_3294_),
    .A2(_3464_),
    .A3(_3335_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7188_ (.I(_3549_),
    .Z(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7189_ (.I0(_3523_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][0] ),
    .S(_3550_),
    .Z(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7190_ (.I(_3551_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7191_ (.I0(_3527_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][1] ),
    .S(_3550_),
    .Z(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7192_ (.I(_3552_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7193_ (.I(_3549_),
    .Z(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7194_ (.I0(_3529_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][2] ),
    .S(_3553_),
    .Z(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7195_ (.I(_3554_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7196_ (.I(_3308_),
    .Z(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7197_ (.A1(_3555_),
    .A2(_3550_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7198_ (.A1(_2206_),
    .A2(_3550_),
    .B(_3556_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7199_ (.I0(_3533_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][4] ),
    .S(_3553_),
    .Z(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7200_ (.I(_3557_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7201_ (.I0(_3508_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][5] ),
    .S(_3553_),
    .Z(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7202_ (.I(_3558_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7203_ (.I0(_3537_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][6] ),
    .S(_3553_),
    .Z(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7204_ (.I(_3559_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7205_ (.I0(_3539_),
    .I1(\mod.Data_Mem.F_M.MRAM[29][7] ),
    .S(_3549_),
    .Z(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7206_ (.I(_3560_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7207_ (.A1(_3270_),
    .A2(_3272_),
    .A3(_3389_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7208_ (.I(_3561_),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7209_ (.I0(_3523_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][0] ),
    .S(_3562_),
    .Z(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7210_ (.I(_3563_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7211_ (.I0(_3527_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][1] ),
    .S(_3562_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7212_ (.I(_3564_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7213_ (.I0(_3529_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][2] ),
    .S(_3562_),
    .Z(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7214_ (.I(_3565_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7215_ (.I0(_3531_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][3] ),
    .S(_3562_),
    .Z(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7216_ (.I(_3566_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7217_ (.I(_3561_),
    .Z(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7218_ (.I0(_3533_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][4] ),
    .S(_3567_),
    .Z(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7219_ (.I(_3568_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7220_ (.I(_3252_),
    .Z(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7221_ (.I0(_3569_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][5] ),
    .S(_3567_),
    .Z(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7222_ (.I(_3570_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7223_ (.I0(_3537_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][6] ),
    .S(_3567_),
    .Z(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7224_ (.I(_3571_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7225_ (.I0(_3539_),
    .I1(\mod.Data_Mem.F_M.MRAM[2][7] ),
    .S(_3567_),
    .Z(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7226_ (.I(_3572_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7227_ (.A1(_3230_),
    .A2(_3464_),
    .A3(_3389_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7228_ (.I(_3573_),
    .Z(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7229_ (.I0(_3523_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][0] ),
    .S(_3574_),
    .Z(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7230_ (.I(_3575_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7231_ (.I0(_3527_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][1] ),
    .S(_3574_),
    .Z(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7232_ (.I(_3576_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7233_ (.I0(_3529_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][2] ),
    .S(_3574_),
    .Z(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7234_ (.I(_3577_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7235_ (.I0(_3531_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][3] ),
    .S(_3574_),
    .Z(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7236_ (.I(_3578_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7237_ (.I(_3573_),
    .Z(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7238_ (.I0(_3533_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][4] ),
    .S(_3579_),
    .Z(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7239_ (.I(_3580_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7240_ (.I0(_3569_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][5] ),
    .S(_3579_),
    .Z(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7241_ (.I(_3581_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7242_ (.I0(_3537_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][6] ),
    .S(_3579_),
    .Z(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7243_ (.I(_3582_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7244_ (.I0(_3539_),
    .I1(\mod.Data_Mem.F_M.MRAM[30][7] ),
    .S(_3579_),
    .Z(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7245_ (.I(_3583_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7246_ (.A1(_3294_),
    .A2(_3464_),
    .A3(_3296_),
    .Z(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7247_ (.I(_3584_),
    .Z(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7248_ (.I0(\mod.Data_Mem.F_M.MRAM[31][0] ),
    .I1(_3293_),
    .S(_3585_),
    .Z(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7249_ (.I(_3586_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7250_ (.I0(_1634_),
    .I1(_3303_),
    .S(_3585_),
    .Z(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7251_ (.I(_3587_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7252_ (.I0(\mod.Data_Mem.F_M.MRAM[31][2] ),
    .I1(_3306_),
    .S(_3585_),
    .Z(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7253_ (.I(_3588_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7254_ (.I0(\mod.Data_Mem.F_M.MRAM[31][3] ),
    .I1(_3555_),
    .S(_3585_),
    .Z(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7255_ (.I(_3589_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7256_ (.I(_3584_),
    .Z(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7257_ (.I0(\mod.Data_Mem.F_M.MRAM[31][4] ),
    .I1(_3312_),
    .S(_3590_),
    .Z(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7258_ (.I(_3591_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7259_ (.I0(\mod.Data_Mem.F_M.MRAM[31][5] ),
    .I1(_3316_),
    .S(_3590_),
    .Z(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7260_ (.I(_3592_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7261_ (.I0(\mod.Data_Mem.F_M.MRAM[31][6] ),
    .I1(_3319_),
    .S(_3590_),
    .Z(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7262_ (.I(_3593_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7263_ (.I0(\mod.Data_Mem.F_M.MRAM[31][7] ),
    .I1(_3322_),
    .S(_3590_),
    .Z(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7264_ (.I(_3594_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7265_ (.I(\mod.Data_Mem.F_M.MRAM[5][0] ),
    .Z(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7266_ (.I(_3595_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7267_ (.I(\mod.Data_Mem.F_M.MRAM[5][1] ),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7268_ (.I(_3596_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7269_ (.I(\mod.Data_Mem.F_M.MRAM[5][2] ),
    .Z(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7270_ (.I(_3597_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7271_ (.I(\mod.Data_Mem.F_M.MRAM[5][3] ),
    .Z(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7272_ (.I(_3598_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7273_ (.I(\mod.Data_Mem.F_M.MRAM[5][4] ),
    .Z(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7274_ (.I(_3599_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7275_ (.I(\mod.Data_Mem.F_M.MRAM[5][5] ),
    .Z(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7276_ (.I(_3600_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7277_ (.I(\mod.Data_Mem.F_M.MRAM[5][6] ),
    .Z(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7278_ (.I(_3601_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7279_ (.I(\mod.Data_Mem.F_M.MRAM[5][7] ),
    .Z(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7280_ (.I(_3602_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7281_ (.I(_3292_),
    .Z(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7282_ (.I(_3297_),
    .Z(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7283_ (.A1(_3232_),
    .A2(_3332_),
    .A3(_3604_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7284_ (.I(_3605_),
    .Z(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7285_ (.I0(_3603_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][0] ),
    .S(_3606_),
    .Z(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7286_ (.I(_3607_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7287_ (.I(_3605_),
    .Z(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7288_ (.I(_3608_),
    .Z(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7289_ (.I(_3302_),
    .Z(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7290_ (.A1(_3610_),
    .A2(_3609_),
    .ZN(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7291_ (.A1(_1719_),
    .A2(_3609_),
    .B(_3611_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7292_ (.I(_3305_),
    .Z(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7293_ (.A1(_3612_),
    .A2(_3606_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7294_ (.A1(_1775_),
    .A2(_3609_),
    .B(_3613_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7295_ (.A1(_3555_),
    .A2(_3606_),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7296_ (.A1(_1855_),
    .A2(_3609_),
    .B(_3614_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7297_ (.I(_3311_),
    .Z(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7298_ (.I0(_3615_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][4] ),
    .S(_3606_),
    .Z(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7299_ (.I(_3616_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7300_ (.I0(_3569_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][5] ),
    .S(_3608_),
    .Z(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7301_ (.I(_3617_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7302_ (.I(_3318_),
    .Z(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7303_ (.I0(_3618_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][6] ),
    .S(_3608_),
    .Z(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7304_ (.I(_3619_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7305_ (.I(_3321_),
    .Z(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7306_ (.I0(_3620_),
    .I1(\mod.Data_Mem.F_M.MRAM[768][7] ),
    .S(_3608_),
    .Z(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7307_ (.I(_3621_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7308_ (.A1(_3332_),
    .A2(_3604_),
    .A3(_3446_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7309_ (.I(_3622_),
    .Z(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7310_ (.I0(_3603_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][0] ),
    .S(_3623_),
    .Z(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7311_ (.I(_3624_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7312_ (.I(_3622_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7313_ (.I(_3625_),
    .Z(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7314_ (.A1(_3610_),
    .A2(_3626_),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7315_ (.A1(_1713_),
    .A2(_3626_),
    .B(_3627_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7316_ (.A1(_3612_),
    .A2(_3623_),
    .ZN(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7317_ (.A1(_1770_),
    .A2(_3626_),
    .B(_3628_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7318_ (.A1(_3555_),
    .A2(_3623_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7319_ (.A1(_1851_),
    .A2(_3626_),
    .B(_3629_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7320_ (.I0(_3615_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][4] ),
    .S(_3623_),
    .Z(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7321_ (.I(_3630_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7322_ (.I0(_3569_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][5] ),
    .S(_3625_),
    .Z(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7323_ (.I(_3631_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7324_ (.I0(_3618_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][6] ),
    .S(_3625_),
    .Z(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7325_ (.I(_3632_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7326_ (.I0(_3620_),
    .I1(\mod.Data_Mem.F_M.MRAM[770][7] ),
    .S(_3625_),
    .Z(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7327_ (.I(_3633_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7328_ (.I(_3297_),
    .Z(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7329_ (.A1(_3272_),
    .A2(_3296_),
    .A3(_3634_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7330_ (.I(_3635_),
    .Z(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7331_ (.I0(_3603_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][0] ),
    .S(_3636_),
    .Z(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7332_ (.I(_3637_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7333_ (.I(_3302_),
    .Z(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7334_ (.I0(_3638_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][1] ),
    .S(_3636_),
    .Z(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7335_ (.I(_3639_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7336_ (.I(_3305_),
    .Z(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7337_ (.I0(_3640_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][2] ),
    .S(_3636_),
    .Z(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7338_ (.I(_3641_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7339_ (.I0(_3531_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][3] ),
    .S(_3636_),
    .Z(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7340_ (.I(_3642_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7341_ (.I(_3635_),
    .Z(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7342_ (.I0(_3615_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][4] ),
    .S(_3643_),
    .Z(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7343_ (.I(_3644_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7344_ (.I(_3315_),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7345_ (.I0(_3645_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][5] ),
    .S(_3643_),
    .Z(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7346_ (.I(_3646_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7347_ (.I0(_3618_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][6] ),
    .S(_3643_),
    .Z(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7348_ (.I(_3647_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7349_ (.I0(_3620_),
    .I1(\mod.Data_Mem.F_M.MRAM[771][7] ),
    .S(_3643_),
    .Z(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7350_ (.I(_3648_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7351_ (.I(\mod.Data_Mem.F_M.MRAM[772][0] ),
    .Z(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7352_ (.I(_3649_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7353_ (.I(\mod.Data_Mem.F_M.MRAM[772][1] ),
    .Z(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7354_ (.I(_3650_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7355_ (.I(\mod.Data_Mem.F_M.MRAM[772][2] ),
    .Z(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7356_ (.I(_3651_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7357_ (.I(\mod.Data_Mem.F_M.MRAM[772][3] ),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7358_ (.I(_3652_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7359_ (.I(\mod.Data_Mem.F_M.MRAM[772][4] ),
    .Z(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7360_ (.I(_3653_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7361_ (.I(\mod.Data_Mem.F_M.MRAM[772][5] ),
    .Z(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7362_ (.I(_3654_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7363_ (.I(\mod.Data_Mem.F_M.MRAM[772][6] ),
    .Z(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7364_ (.I(_3655_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7365_ (.I(\mod.Data_Mem.F_M.MRAM[772][7] ),
    .Z(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7366_ (.I(_3656_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7367_ (.I(\mod.Data_Mem.F_M.MRAM[773][0] ),
    .Z(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7368_ (.I(_3657_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7369_ (.I(\mod.Data_Mem.F_M.MRAM[773][1] ),
    .Z(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7370_ (.I(_3658_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7371_ (.I(\mod.Data_Mem.F_M.MRAM[773][2] ),
    .Z(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7372_ (.I(_3659_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7373_ (.I(\mod.Data_Mem.F_M.MRAM[773][3] ),
    .Z(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7374_ (.I(_3660_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7375_ (.I(\mod.Data_Mem.F_M.MRAM[773][4] ),
    .Z(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7376_ (.I(_3661_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7377_ (.I(\mod.Data_Mem.F_M.MRAM[773][5] ),
    .Z(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7378_ (.I(_3662_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7379_ (.I(\mod.Data_Mem.F_M.MRAM[773][6] ),
    .Z(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7380_ (.I(_3663_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7381_ (.I(\mod.Data_Mem.F_M.MRAM[773][7] ),
    .Z(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7382_ (.I(_3664_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7383_ (.I(\mod.Data_Mem.F_M.MRAM[774][0] ),
    .Z(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7384_ (.I(_3665_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7385_ (.I(\mod.Data_Mem.F_M.MRAM[774][1] ),
    .Z(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7386_ (.I(_3666_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7387_ (.I(\mod.Data_Mem.F_M.MRAM[774][2] ),
    .Z(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7388_ (.I(_3667_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7389_ (.I(\mod.Data_Mem.F_M.MRAM[774][3] ),
    .Z(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7390_ (.I(_3668_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7391_ (.I(\mod.Data_Mem.F_M.MRAM[774][4] ),
    .Z(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7392_ (.I(_3669_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7393_ (.I(\mod.Data_Mem.F_M.MRAM[774][5] ),
    .Z(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7394_ (.I(_3670_),
    .Z(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7395_ (.I(\mod.Data_Mem.F_M.MRAM[774][6] ),
    .Z(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7396_ (.I(_3671_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7397_ (.I(\mod.Data_Mem.F_M.MRAM[774][7] ),
    .Z(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7398_ (.I(_3672_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7399_ (.I(\mod.Data_Mem.F_M.MRAM[775][0] ),
    .Z(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7400_ (.I(_3673_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7401_ (.I(\mod.Data_Mem.F_M.MRAM[775][1] ),
    .Z(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7402_ (.I(_3674_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7403_ (.I(\mod.Data_Mem.F_M.MRAM[775][2] ),
    .Z(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7404_ (.I(_3675_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7405_ (.I(\mod.Data_Mem.F_M.MRAM[775][3] ),
    .Z(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7406_ (.I(_3676_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7407_ (.I(\mod.Data_Mem.F_M.MRAM[775][4] ),
    .Z(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7408_ (.I(_3677_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7409_ (.I(\mod.Data_Mem.F_M.MRAM[775][5] ),
    .Z(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7410_ (.I(_3678_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7411_ (.I(\mod.Data_Mem.F_M.MRAM[775][6] ),
    .Z(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7412_ (.I(_3679_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7413_ (.I(\mod.Data_Mem.F_M.MRAM[775][7] ),
    .Z(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7414_ (.I(_3680_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7415_ (.I(\mod.Data_Mem.F_M.MRAM[776][0] ),
    .Z(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7416_ (.I(_3681_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7417_ (.I(\mod.Data_Mem.F_M.MRAM[776][1] ),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7418_ (.I(_3682_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7419_ (.I(\mod.Data_Mem.F_M.MRAM[776][2] ),
    .Z(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7420_ (.I(_3683_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7421_ (.I(\mod.Data_Mem.F_M.MRAM[776][3] ),
    .Z(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7422_ (.I(_3684_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7423_ (.I(\mod.Data_Mem.F_M.MRAM[776][4] ),
    .Z(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7424_ (.I(_3685_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7425_ (.I(\mod.Data_Mem.F_M.MRAM[776][5] ),
    .Z(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7426_ (.I(_3686_),
    .Z(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7427_ (.I(\mod.Data_Mem.F_M.MRAM[776][6] ),
    .Z(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7428_ (.I(_3687_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7429_ (.I(\mod.Data_Mem.F_M.MRAM[776][7] ),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7430_ (.I(_3688_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7431_ (.I(\mod.Data_Mem.F_M.MRAM[777][0] ),
    .Z(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7432_ (.I(_3689_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7433_ (.I(\mod.Data_Mem.F_M.MRAM[777][1] ),
    .Z(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7434_ (.I(_3690_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7435_ (.I(\mod.Data_Mem.F_M.MRAM[777][2] ),
    .Z(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7436_ (.I(_3691_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7437_ (.I(\mod.Data_Mem.F_M.MRAM[777][3] ),
    .Z(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7438_ (.I(_3692_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7439_ (.I(\mod.Data_Mem.F_M.MRAM[777][4] ),
    .Z(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7440_ (.I(_3693_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7441_ (.I(\mod.Data_Mem.F_M.MRAM[777][5] ),
    .Z(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7442_ (.I(_3694_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7443_ (.I(\mod.Data_Mem.F_M.MRAM[777][6] ),
    .Z(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7444_ (.I(_3695_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7445_ (.I(\mod.Data_Mem.F_M.MRAM[777][7] ),
    .Z(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7446_ (.I(_3696_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7447_ (.I(\mod.Data_Mem.F_M.MRAM[778][0] ),
    .Z(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7448_ (.I(_3697_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7449_ (.I(\mod.Data_Mem.F_M.MRAM[778][1] ),
    .Z(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7450_ (.I(_3698_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7451_ (.I(\mod.Data_Mem.F_M.MRAM[778][2] ),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7452_ (.I(_3699_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7453_ (.I(\mod.Data_Mem.F_M.MRAM[778][3] ),
    .Z(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7454_ (.I(_3700_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7455_ (.I(\mod.Data_Mem.F_M.MRAM[778][4] ),
    .Z(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7456_ (.I(_3701_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7457_ (.I(\mod.Data_Mem.F_M.MRAM[778][5] ),
    .Z(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7458_ (.I(_3702_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7459_ (.I(\mod.Data_Mem.F_M.MRAM[778][6] ),
    .Z(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7460_ (.I(_3703_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7461_ (.I(\mod.Data_Mem.F_M.MRAM[778][7] ),
    .Z(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7462_ (.I(_3704_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7463_ (.I(_3297_),
    .Z(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7464_ (.A1(_3269_),
    .A2(_3705_),
    .A3(_3374_),
    .ZN(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7465_ (.I(_3706_),
    .Z(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7466_ (.I0(_3603_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][0] ),
    .S(_3707_),
    .Z(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7467_ (.I(_3708_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7468_ (.I0(_3638_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][1] ),
    .S(_3707_),
    .Z(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7469_ (.I(_3709_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7470_ (.I0(_3640_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][2] ),
    .S(_3707_),
    .Z(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7471_ (.I(_3710_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7472_ (.I(_3308_),
    .Z(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7473_ (.I0(_3711_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][3] ),
    .S(_3707_),
    .Z(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7474_ (.I(_3712_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7475_ (.I(_3706_),
    .Z(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7476_ (.I0(_3615_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][4] ),
    .S(_3713_),
    .Z(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7477_ (.I(_3714_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7478_ (.I0(_3645_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][5] ),
    .S(_3713_),
    .Z(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7479_ (.I(_3715_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7480_ (.I0(_3618_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][6] ),
    .S(_3713_),
    .Z(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7481_ (.I(_3716_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7482_ (.I0(_3620_),
    .I1(\mod.Data_Mem.F_M.MRAM[780][7] ),
    .S(_3713_),
    .Z(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7483_ (.I(_3717_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7484_ (.I(_3292_),
    .Z(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7485_ (.A1(_3634_),
    .A2(_3371_),
    .A3(_3387_),
    .ZN(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7486_ (.I(_3719_),
    .Z(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7487_ (.I0(_3718_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][0] ),
    .S(_3720_),
    .Z(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7488_ (.I(_3721_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7489_ (.I0(_3638_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][1] ),
    .S(_3720_),
    .Z(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7490_ (.I(_3722_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7491_ (.I0(_3640_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][2] ),
    .S(_3720_),
    .Z(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7492_ (.I(_3723_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7493_ (.I0(_3711_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][3] ),
    .S(_3720_),
    .Z(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7494_ (.I(_3724_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7495_ (.I(_3311_),
    .Z(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7496_ (.I(_3719_),
    .Z(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7497_ (.I0(_3725_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][4] ),
    .S(_3726_),
    .Z(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7498_ (.I(_3727_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7499_ (.I0(_3645_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][5] ),
    .S(_3726_),
    .Z(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7500_ (.I(_3728_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7501_ (.I(_3318_),
    .Z(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7502_ (.I0(_3729_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][6] ),
    .S(_3726_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7503_ (.I(_3730_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7504_ (.I(_3321_),
    .Z(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7505_ (.I0(_3731_),
    .I1(\mod.Data_Mem.F_M.MRAM[781][7] ),
    .S(_3726_),
    .Z(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7506_ (.I(_3732_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7507_ (.A1(_3634_),
    .A2(_3387_),
    .A3(_3389_),
    .ZN(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7508_ (.I(_3733_),
    .Z(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7509_ (.I0(_3718_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][0] ),
    .S(_3734_),
    .Z(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7510_ (.I(_3735_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7511_ (.I0(_3638_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][1] ),
    .S(_3734_),
    .Z(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7512_ (.I(_3736_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7513_ (.I0(_3640_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][2] ),
    .S(_3734_),
    .Z(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7514_ (.I(_3737_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7515_ (.I0(_3711_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][3] ),
    .S(_3734_),
    .Z(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7516_ (.I(_3738_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7517_ (.I(_3733_),
    .Z(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7518_ (.I0(_3725_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][4] ),
    .S(_3739_),
    .Z(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7519_ (.I(_3740_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7520_ (.I0(_3645_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][5] ),
    .S(_3739_),
    .Z(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7521_ (.I(_3741_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7522_ (.I0(_3729_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][6] ),
    .S(_3739_),
    .Z(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7523_ (.I(_3742_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7524_ (.I0(_3731_),
    .I1(\mod.Data_Mem.F_M.MRAM[782][7] ),
    .S(_3739_),
    .Z(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7525_ (.I(_3743_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7526_ (.A1(_3407_),
    .A2(_3705_),
    .A3(_3387_),
    .ZN(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7527_ (.I(_3744_),
    .Z(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7528_ (.I0(_3718_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][0] ),
    .S(_3745_),
    .Z(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7529_ (.I(_3746_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7530_ (.I(_3302_),
    .Z(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7531_ (.I0(_3747_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][1] ),
    .S(_3745_),
    .Z(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7532_ (.I(_3748_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7533_ (.I(_3305_),
    .Z(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7534_ (.I0(_3749_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][2] ),
    .S(_3745_),
    .Z(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7535_ (.I(_3750_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7536_ (.I0(_3711_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][3] ),
    .S(_3745_),
    .Z(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7537_ (.I(_3751_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7538_ (.I(_3744_),
    .Z(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7539_ (.I0(_3725_),
    .I1(_1902_),
    .S(_3752_),
    .Z(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7540_ (.I(_3753_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7541_ (.I(_3315_),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7542_ (.I0(_3754_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][5] ),
    .S(_3752_),
    .Z(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7543_ (.I(_3755_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7544_ (.I0(_3729_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][6] ),
    .S(_3752_),
    .Z(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7545_ (.I(_3756_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7546_ (.I0(_3731_),
    .I1(\mod.Data_Mem.F_M.MRAM[783][7] ),
    .S(_3752_),
    .Z(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7547_ (.I(_3757_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7548_ (.I(_3420_),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7549_ (.A1(_3232_),
    .A2(_3298_),
    .A3(_3758_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7550_ (.I(_3759_),
    .Z(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7551_ (.I0(_3718_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][0] ),
    .S(_3760_),
    .Z(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7552_ (.I(_3761_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7553_ (.I(_3759_),
    .Z(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7554_ (.A1(_3610_),
    .A2(_3762_),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7555_ (.A1(_1683_),
    .A2(_3762_),
    .B(_3763_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7556_ (.A1(_3612_),
    .A2(_3762_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7557_ (.A1(_1797_),
    .A2(_3762_),
    .B(_3764_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7558_ (.I(_3308_),
    .Z(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7559_ (.I0(_3765_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][3] ),
    .S(_3760_),
    .Z(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7560_ (.I(_3766_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7561_ (.I0(_3725_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][4] ),
    .S(_3760_),
    .Z(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7562_ (.I(_3767_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7563_ (.I0(_3754_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][5] ),
    .S(_3760_),
    .Z(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7564_ (.I(_3768_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7565_ (.I0(_3729_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][6] ),
    .S(_3759_),
    .Z(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7566_ (.I(_3769_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7567_ (.I0(_3731_),
    .I1(\mod.Data_Mem.F_M.MRAM[784][7] ),
    .S(_3759_),
    .Z(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7568_ (.I(_3770_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7569_ (.I(_3292_),
    .Z(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7570_ (.A1(_3705_),
    .A2(_3335_),
    .A3(_3758_),
    .ZN(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7571_ (.I(_3772_),
    .Z(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7572_ (.I0(_3771_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][0] ),
    .S(_3773_),
    .Z(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7573_ (.I(_3774_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7574_ (.I0(_3747_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][1] ),
    .S(_3773_),
    .Z(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7575_ (.I(_3775_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7576_ (.I0(_3749_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][2] ),
    .S(_3773_),
    .Z(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7577_ (.I(_3776_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7578_ (.I0(_3765_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][3] ),
    .S(_3773_),
    .Z(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7579_ (.I(_3777_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7580_ (.I(_3311_),
    .Z(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7581_ (.I(_3772_),
    .Z(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7582_ (.I0(_3778_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][4] ),
    .S(_3779_),
    .Z(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7583_ (.I(_3780_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7584_ (.I0(_3754_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][5] ),
    .S(_3779_),
    .Z(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7585_ (.I(_3781_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7586_ (.I(_3318_),
    .Z(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7587_ (.I0(_3782_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][6] ),
    .S(_3779_),
    .Z(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7588_ (.I(_3783_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7589_ (.I(_3321_),
    .Z(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7590_ (.I0(_3784_),
    .I1(\mod.Data_Mem.F_M.MRAM[785][7] ),
    .S(_3779_),
    .Z(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7591_ (.I(_3785_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7592_ (.A1(_3604_),
    .A2(_3446_),
    .A3(_3758_),
    .ZN(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7593_ (.I(_3786_),
    .Z(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7594_ (.I0(_3771_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][0] ),
    .S(_3787_),
    .Z(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7595_ (.I(_3788_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7596_ (.I(_3786_),
    .Z(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7597_ (.A1(_3610_),
    .A2(_3789_),
    .ZN(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7598_ (.A1(_1686_),
    .A2(_3789_),
    .B(_3790_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7599_ (.A1(_3612_),
    .A2(_3789_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7600_ (.A1(_1793_),
    .A2(_3789_),
    .B(_3791_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7601_ (.I0(_3765_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][3] ),
    .S(_3787_),
    .Z(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7602_ (.I(_3792_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7603_ (.I0(_3778_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][4] ),
    .S(_3787_),
    .Z(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7604_ (.I(_3793_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7605_ (.I0(_3754_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][5] ),
    .S(_3787_),
    .Z(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7606_ (.I(_3794_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7607_ (.I0(_3782_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][6] ),
    .S(_3786_),
    .Z(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7608_ (.I(_3795_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7609_ (.I0(_3784_),
    .I1(\mod.Data_Mem.F_M.MRAM[786][7] ),
    .S(_3786_),
    .Z(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7610_ (.I(_3796_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7611_ (.A1(_3296_),
    .A2(_3604_),
    .A3(_3758_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7612_ (.I(_3797_),
    .Z(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7613_ (.I0(_3771_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][0] ),
    .S(_3798_),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7614_ (.I(_3799_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7615_ (.I0(_3747_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][1] ),
    .S(_3798_),
    .Z(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7616_ (.I(_3800_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7617_ (.I(_3797_),
    .Z(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7618_ (.I0(_3749_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][2] ),
    .S(_3801_),
    .Z(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7619_ (.I(_3802_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7620_ (.I0(_3765_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][3] ),
    .S(_3801_),
    .Z(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7621_ (.I(_3803_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7622_ (.I(_3801_),
    .Z(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7623_ (.A1(_3312_),
    .A2(_3804_),
    .ZN(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7624_ (.A1(_1922_),
    .A2(_3804_),
    .B(_3805_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7625_ (.I(_3315_),
    .Z(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7626_ (.I0(_3806_),
    .I1(\mod.Data_Mem.F_M.MRAM[787][5] ),
    .S(_3801_),
    .Z(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7627_ (.I(_3807_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7628_ (.A1(_3319_),
    .A2(_3798_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7629_ (.A1(_2009_),
    .A2(_3804_),
    .B(_3808_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7630_ (.A1(_3322_),
    .A2(_3798_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7631_ (.A1(_2043_),
    .A2(_3804_),
    .B(_3809_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7632_ (.I(\mod.Data_Mem.F_M.MRAM[788][0] ),
    .Z(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7633_ (.I(_3810_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7634_ (.I(\mod.Data_Mem.F_M.MRAM[788][1] ),
    .Z(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7635_ (.I(_3811_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7636_ (.I(\mod.Data_Mem.F_M.MRAM[788][2] ),
    .Z(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7637_ (.I(_3812_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7638_ (.I(\mod.Data_Mem.F_M.MRAM[788][3] ),
    .Z(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7639_ (.I(_3813_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7640_ (.I(\mod.Data_Mem.F_M.MRAM[788][4] ),
    .Z(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7641_ (.I(_3814_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7642_ (.I(\mod.Data_Mem.F_M.MRAM[788][5] ),
    .Z(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7643_ (.I(_3815_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7644_ (.I(\mod.Data_Mem.F_M.MRAM[788][6] ),
    .Z(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7645_ (.I(_3816_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7646_ (.I(\mod.Data_Mem.F_M.MRAM[788][7] ),
    .Z(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7647_ (.I(_3817_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7648_ (.I(\mod.Data_Mem.F_M.MRAM[790][0] ),
    .Z(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7649_ (.I(_3818_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7650_ (.I(\mod.Data_Mem.F_M.MRAM[790][1] ),
    .Z(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7651_ (.I(_3819_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7652_ (.I(\mod.Data_Mem.F_M.MRAM[790][2] ),
    .Z(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7653_ (.I(_3820_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7654_ (.I(\mod.Data_Mem.F_M.MRAM[790][3] ),
    .Z(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7655_ (.I(_3821_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7656_ (.I(\mod.Data_Mem.F_M.MRAM[790][4] ),
    .Z(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7657_ (.I(_3822_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7658_ (.I(\mod.Data_Mem.F_M.MRAM[790][5] ),
    .Z(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7659_ (.I(_3823_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7660_ (.I(\mod.Data_Mem.F_M.MRAM[790][6] ),
    .Z(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7661_ (.I(_3824_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7662_ (.I(\mod.Data_Mem.F_M.MRAM[790][7] ),
    .Z(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7663_ (.I(_3825_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7664_ (.I(\mod.Data_Mem.F_M.MRAM[791][0] ),
    .Z(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7665_ (.I(_3826_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7666_ (.I(\mod.Data_Mem.F_M.MRAM[791][1] ),
    .Z(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7667_ (.I(_3827_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7668_ (.I(\mod.Data_Mem.F_M.MRAM[791][2] ),
    .Z(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7669_ (.I(_3828_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7670_ (.I(\mod.Data_Mem.F_M.MRAM[791][3] ),
    .Z(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7671_ (.I(_3829_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7672_ (.I(\mod.Data_Mem.F_M.MRAM[791][4] ),
    .Z(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7673_ (.I(_3830_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7674_ (.I(\mod.Data_Mem.F_M.MRAM[791][5] ),
    .Z(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7675_ (.I(_3831_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7676_ (.I(\mod.Data_Mem.F_M.MRAM[791][6] ),
    .Z(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7677_ (.I(_3832_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7678_ (.I(\mod.Data_Mem.F_M.MRAM[791][7] ),
    .Z(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7679_ (.I(_3833_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7680_ (.I(\mod.Data_Mem.F_M.MRAM[792][0] ),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7681_ (.I(_3834_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7682_ (.I(\mod.Data_Mem.F_M.MRAM[792][1] ),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7683_ (.I(_3835_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7684_ (.I(\mod.Data_Mem.F_M.MRAM[792][2] ),
    .Z(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7685_ (.I(_3836_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7686_ (.I(\mod.Data_Mem.F_M.MRAM[792][3] ),
    .Z(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7687_ (.I(_3837_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7688_ (.I(\mod.Data_Mem.F_M.MRAM[792][4] ),
    .Z(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7689_ (.I(_3838_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7690_ (.I(\mod.Data_Mem.F_M.MRAM[792][5] ),
    .Z(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7691_ (.I(_3839_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7692_ (.I(\mod.Data_Mem.F_M.MRAM[792][6] ),
    .Z(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7693_ (.I(_3840_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7694_ (.I(\mod.Data_Mem.F_M.MRAM[792][7] ),
    .Z(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7695_ (.I(_3841_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7696_ (.I(\mod.Data_Mem.F_M.MRAM[793][0] ),
    .Z(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7697_ (.I(_3842_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7698_ (.I(\mod.Data_Mem.F_M.MRAM[793][1] ),
    .Z(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7699_ (.I(_3843_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7700_ (.I(\mod.Data_Mem.F_M.MRAM[793][2] ),
    .Z(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7701_ (.I(_3844_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7702_ (.I(\mod.Data_Mem.F_M.MRAM[793][3] ),
    .Z(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7703_ (.I(_3845_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7704_ (.I(\mod.Data_Mem.F_M.MRAM[793][4] ),
    .Z(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7705_ (.I(_3846_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7706_ (.I(\mod.Data_Mem.F_M.MRAM[793][5] ),
    .Z(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7707_ (.I(_3847_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7708_ (.I(\mod.Data_Mem.F_M.MRAM[793][6] ),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7709_ (.I(_3848_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7710_ (.I(\mod.Data_Mem.F_M.MRAM[793][7] ),
    .Z(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7711_ (.I(_3849_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7712_ (.I(\mod.Data_Mem.F_M.MRAM[794][0] ),
    .Z(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7713_ (.I(_3850_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7714_ (.I(\mod.Data_Mem.F_M.MRAM[794][1] ),
    .Z(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7715_ (.I(_3851_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7716_ (.I(\mod.Data_Mem.F_M.MRAM[794][2] ),
    .Z(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7717_ (.I(_3852_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7718_ (.I(\mod.Data_Mem.F_M.MRAM[794][3] ),
    .Z(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7719_ (.I(_3853_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7720_ (.I(\mod.Data_Mem.F_M.MRAM[794][4] ),
    .Z(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7721_ (.I(_3854_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7722_ (.I(\mod.Data_Mem.F_M.MRAM[794][5] ),
    .Z(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7723_ (.I(_3855_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7724_ (.I(\mod.Data_Mem.F_M.MRAM[794][6] ),
    .Z(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7725_ (.I(_3856_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7726_ (.I(\mod.Data_Mem.F_M.MRAM[794][7] ),
    .Z(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7727_ (.I(_3857_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7728_ (.I(\mod.Data_Mem.F_M.MRAM[795][0] ),
    .Z(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7729_ (.I(_3858_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7730_ (.I(\mod.Data_Mem.F_M.MRAM[795][1] ),
    .Z(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7731_ (.I(_3859_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7732_ (.I(\mod.Data_Mem.F_M.MRAM[795][2] ),
    .Z(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7733_ (.I(_3860_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7734_ (.I(\mod.Data_Mem.F_M.MRAM[795][3] ),
    .Z(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7735_ (.I(_3861_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7736_ (.I(\mod.Data_Mem.F_M.MRAM[795][4] ),
    .Z(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7737_ (.I(_3862_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7738_ (.I(\mod.Data_Mem.F_M.MRAM[795][5] ),
    .Z(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7739_ (.I(_3863_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7740_ (.I(\mod.Data_Mem.F_M.MRAM[795][6] ),
    .Z(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7741_ (.I(_3864_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7742_ (.I(\mod.Data_Mem.F_M.MRAM[795][7] ),
    .Z(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7743_ (.I(_3865_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7744_ (.A1(_3230_),
    .A2(_3232_),
    .A3(_3634_),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7745_ (.I(_3866_),
    .Z(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7746_ (.I0(_3771_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][0] ),
    .S(_3867_),
    .Z(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7747_ (.I(_3868_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7748_ (.I0(_3747_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][1] ),
    .S(_3867_),
    .Z(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7749_ (.I(_3869_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7750_ (.I0(_3749_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][2] ),
    .S(_3867_),
    .Z(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7751_ (.I(_3870_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7752_ (.I0(_3309_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][3] ),
    .S(_3867_),
    .Z(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7753_ (.I(_3871_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7754_ (.I(_3866_),
    .Z(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7755_ (.I0(_3778_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][4] ),
    .S(_3872_),
    .Z(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7756_ (.I(_3873_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7757_ (.I0(_3806_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][5] ),
    .S(_3872_),
    .Z(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7758_ (.I(_3874_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7759_ (.I0(_3782_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][6] ),
    .S(_3872_),
    .Z(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7760_ (.I(_3875_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7761_ (.I0(_3784_),
    .I1(\mod.Data_Mem.F_M.MRAM[796][7] ),
    .S(_3872_),
    .Z(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7762_ (.I(_3876_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7763_ (.A1(_3230_),
    .A2(_3705_),
    .A3(_3371_),
    .ZN(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7764_ (.I(_3877_),
    .Z(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7765_ (.I0(_3293_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][0] ),
    .S(_3878_),
    .Z(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7766_ (.I(_3879_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7767_ (.I0(_3303_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][1] ),
    .S(_3878_),
    .Z(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7768_ (.I(_3880_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7769_ (.I0(_3306_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][2] ),
    .S(_3878_),
    .Z(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7770_ (.I(_3881_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7771_ (.I0(_3309_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][3] ),
    .S(_3878_),
    .Z(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7772_ (.I(_3882_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7773_ (.I(_3877_),
    .Z(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7774_ (.I0(_3778_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][4] ),
    .S(_3883_),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7775_ (.I(_3884_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7776_ (.I0(_3806_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][5] ),
    .S(_3883_),
    .Z(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7777_ (.I(_3885_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7778_ (.I0(_3782_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][6] ),
    .S(_3883_),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7779_ (.I(_3886_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7780_ (.I0(_3784_),
    .I1(\mod.Data_Mem.F_M.MRAM[797][7] ),
    .S(_3883_),
    .Z(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7781_ (.I(_3887_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7782_ (.A1(_3294_),
    .A2(_3298_),
    .A3(_3446_),
    .ZN(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7783_ (.I(_3888_),
    .Z(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7784_ (.I0(_3293_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][0] ),
    .S(_3889_),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7785_ (.I(_3890_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7786_ (.I0(_3303_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][1] ),
    .S(_3889_),
    .Z(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7787_ (.I(_3891_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7788_ (.I0(_3306_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][2] ),
    .S(_3889_),
    .Z(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7789_ (.I(_3892_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7790_ (.I0(_3309_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][3] ),
    .S(_3889_),
    .Z(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7791_ (.I(_3893_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7792_ (.I(_3888_),
    .Z(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7793_ (.I0(_3312_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][4] ),
    .S(_3894_),
    .Z(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7794_ (.I(_3895_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7795_ (.I0(_3806_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][5] ),
    .S(_3894_),
    .Z(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7796_ (.I(_3896_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7797_ (.I0(_3319_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][6] ),
    .S(_3894_),
    .Z(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7798_ (.I(_3897_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7799_ (.I0(_3322_),
    .I1(\mod.Data_Mem.F_M.MRAM[798][7] ),
    .S(_3894_),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7800_ (.I(_3898_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7801_ (.I(\mod.Data_Mem.F_M.MRAM[7][0] ),
    .Z(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7802_ (.I(_3899_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7803_ (.I(\mod.Data_Mem.F_M.MRAM[7][1] ),
    .Z(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7804_ (.I(_3900_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7805_ (.I(\mod.Data_Mem.F_M.MRAM[7][2] ),
    .Z(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7806_ (.I(_3901_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7807_ (.I(\mod.Data_Mem.F_M.MRAM[7][3] ),
    .Z(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7808_ (.I(_3902_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7809_ (.I(\mod.Data_Mem.F_M.MRAM[7][4] ),
    .Z(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7810_ (.I(_3903_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7811_ (.I(\mod.Data_Mem.F_M.MRAM[7][5] ),
    .Z(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7812_ (.I(_3904_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7813_ (.I(\mod.Data_Mem.F_M.MRAM[7][6] ),
    .Z(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7814_ (.I(_3905_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7815_ (.I(\mod.Data_Mem.F_M.MRAM[7][7] ),
    .Z(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7816_ (.I(_3906_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7817_ (.I(\mod.I_addr[3] ),
    .Z(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7818_ (.A1(\mod.I_addr[4] ),
    .A2(\mod.I_addr[6] ),
    .A3(\mod.I_addr[5] ),
    .A4(\mod.I_addr[7] ),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7819_ (.A1(\mod.I_addr[0] ),
    .A2(\mod.I_addr[2] ),
    .A3(\mod.I_addr[1] ),
    .ZN(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7820_ (.A1(_3907_),
    .A2(_3908_),
    .A3(_3909_),
    .Z(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7821_ (.I(_3910_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7822_ (.A1(\mod.I_addr[0] ),
    .A2(_3169_),
    .ZN(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7823_ (.A1(_3171_),
    .A2(_3908_),
    .ZN(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7824_ (.A1(_3907_),
    .A2(_3911_),
    .A3(_3912_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7825_ (.A1(_3907_),
    .A2(_3912_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7826_ (.A1(\mod.I_addr[3] ),
    .A2(_3911_),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7827_ (.A1(_3908_),
    .A2(_3913_),
    .Z(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7828_ (.I(_3914_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7829_ (.A1(_3174_),
    .A2(_3909_),
    .B(_3908_),
    .ZN(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7830_ (.I(_3915_),
    .Z(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7831_ (.A1(_0612_),
    .A2(_3175_),
    .B(_3916_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7832_ (.I(_3916_),
    .Z(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7833_ (.A1(_0081_),
    .A2(_3917_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7834_ (.A1(_0080_),
    .A2(_3171_),
    .Z(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7835_ (.A1(_3175_),
    .A2(_3918_),
    .B(_3916_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7836_ (.A1(_3907_),
    .A2(\mod.I_addr[2] ),
    .ZN(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7837_ (.A1(_3913_),
    .A2(_3915_),
    .A3(_3919_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7838_ (.I(_3920_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7839_ (.I(_3169_),
    .ZN(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7840_ (.A1(_0080_),
    .A2(_3171_),
    .B(_3921_),
    .C(_3916_),
    .ZN(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7841_ (.A1(_0610_),
    .A2(_3922_),
    .Z(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7842_ (.I(_3923_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7843_ (.I(\mod.Data_Mem.F_M.MRAM[9][0] ),
    .Z(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7844_ (.I(_3924_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7845_ (.I(\mod.Data_Mem.F_M.MRAM[9][1] ),
    .Z(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7846_ (.I(_3925_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7847_ (.I(\mod.Data_Mem.F_M.MRAM[9][2] ),
    .Z(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7848_ (.I(_3926_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7849_ (.I(\mod.Data_Mem.F_M.MRAM[9][3] ),
    .Z(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7850_ (.I(_3927_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7851_ (.I(\mod.Data_Mem.F_M.MRAM[9][4] ),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7852_ (.I(_3928_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7853_ (.I(\mod.Data_Mem.F_M.MRAM[9][5] ),
    .Z(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7854_ (.I(_3929_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7855_ (.I(\mod.Data_Mem.F_M.MRAM[9][6] ),
    .Z(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7856_ (.I(_3930_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7857_ (.I(\mod.Data_Mem.F_M.MRAM[9][7] ),
    .Z(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7858_ (.I(_3931_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7859_ (.A1(_3913_),
    .A2(_3917_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7860_ (.I(_3917_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7861_ (.A1(_3917_),
    .A2(_3919_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7862_ (.D(_0088_),
    .CLK(net378),
    .Q(\mod.Data_Mem.F_M.MRAM[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7863_ (.D(_0089_),
    .CLK(net382),
    .Q(\mod.Data_Mem.F_M.MRAM[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7864_ (.D(_0090_),
    .CLK(net173),
    .Q(\mod.Data_Mem.F_M.MRAM[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7865_ (.D(_0091_),
    .CLK(net166),
    .Q(\mod.Data_Mem.F_M.MRAM[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7866_ (.D(_0092_),
    .CLK(net167),
    .Q(\mod.Data_Mem.F_M.MRAM[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7867_ (.D(_0093_),
    .CLK(net371),
    .Q(\mod.Data_Mem.F_M.MRAM[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7868_ (.D(_0094_),
    .CLK(net378),
    .Q(\mod.Data_Mem.F_M.MRAM[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7869_ (.D(_0095_),
    .CLK(net320),
    .Q(\mod.Data_Mem.F_M.MRAM[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7870_ (.D(_0096_),
    .CLK(net375),
    .Q(\mod.Data_Mem.F_M.MRAM[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7871_ (.D(_0097_),
    .CLK(net372),
    .Q(\mod.Data_Mem.F_M.MRAM[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7872_ (.D(_0098_),
    .CLK(net320),
    .Q(\mod.Data_Mem.F_M.MRAM[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7873_ (.D(_0099_),
    .CLK(net316),
    .Q(\mod.Data_Mem.F_M.MRAM[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7874_ (.D(_0100_),
    .CLK(net172),
    .Q(\mod.Data_Mem.F_M.MRAM[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7875_ (.D(_0101_),
    .CLK(net156),
    .Q(\mod.Data_Mem.F_M.MRAM[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7876_ (.D(_0102_),
    .CLK(net386),
    .Q(\mod.Data_Mem.F_M.MRAM[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7877_ (.D(_0103_),
    .CLK(net376),
    .Q(\mod.Data_Mem.F_M.MRAM[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7878_ (.D(_0104_),
    .CLK(net372),
    .Q(\mod.Data_Mem.F_M.MRAM[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7879_ (.D(_0105_),
    .CLK(net317),
    .Q(\mod.Data_Mem.F_M.MRAM[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7880_ (.D(_0106_),
    .CLK(net170),
    .Q(\mod.Data_Mem.F_M.MRAM[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7881_ (.D(_0107_),
    .CLK(net321),
    .Q(\mod.Data_Mem.F_M.MRAM[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7882_ (.D(_0108_),
    .CLK(net155),
    .Q(\mod.Data_Mem.F_M.MRAM[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7883_ (.D(_0109_),
    .CLK(net384),
    .Q(\mod.Data_Mem.F_M.MRAM[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7884_ (.D(_0110_),
    .CLK(net376),
    .Q(\mod.Data_Mem.F_M.MRAM[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7885_ (.D(_0111_),
    .CLK(net379),
    .Q(\mod.Data_Mem.F_M.MRAM[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7886_ (.D(_0112_),
    .CLK(net386),
    .Q(\mod.Data_Mem.F_M.MRAM[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7887_ (.D(_0113_),
    .CLK(net157),
    .Q(\mod.Data_Mem.F_M.MRAM[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7888_ (.D(_0114_),
    .CLK(net322),
    .Q(\mod.Data_Mem.F_M.MRAM[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7889_ (.D(_0115_),
    .CLK(net387),
    .Q(\mod.Data_Mem.F_M.MRAM[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7890_ (.D(_0116_),
    .CLK(net170),
    .Q(\mod.Data_Mem.F_M.MRAM[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7891_ (.D(_0117_),
    .CLK(net173),
    .Q(\mod.Data_Mem.F_M.MRAM[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7892_ (.D(_0118_),
    .CLK(net171),
    .Q(\mod.Data_Mem.F_M.MRAM[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7893_ (.D(_0119_),
    .CLK(net383),
    .Q(\mod.Data_Mem.F_M.MRAM[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7894_ (.D(_0120_),
    .CLK(net205),
    .Q(\mod.Data_Mem.F_M.MRAM[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7895_ (.D(_0121_),
    .CLK(net370),
    .Q(\mod.Data_Mem.F_M.MRAM[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7896_ (.D(_0122_),
    .CLK(net369),
    .Q(\mod.Data_Mem.F_M.MRAM[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7897_ (.D(_0123_),
    .CLK(net193),
    .Q(\mod.Data_Mem.F_M.MRAM[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7898_ (.D(_0124_),
    .CLK(net383),
    .Q(\mod.Data_Mem.F_M.MRAM[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7899_ (.D(_0125_),
    .CLK(net197),
    .Q(\mod.Data_Mem.F_M.MRAM[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7900_ (.D(_0126_),
    .CLK(net172),
    .Q(\mod.Data_Mem.F_M.MRAM[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7901_ (.D(_0127_),
    .CLK(net303),
    .Q(\mod.Data_Mem.F_M.MRAM[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7902_ (.D(_0128_),
    .CLK(net307),
    .Q(\mod.Data_Mem.F_M.MRAM[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7903_ (.D(_0129_),
    .CLK(net312),
    .Q(\mod.Data_Mem.F_M.MRAM[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7904_ (.D(_0130_),
    .CLK(net320),
    .Q(\mod.Data_Mem.F_M.MRAM[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7905_ (.D(_0131_),
    .CLK(net307),
    .Q(\mod.Data_Mem.F_M.MRAM[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7906_ (.D(_0132_),
    .CLK(net242),
    .Q(\mod.Data_Mem.F_M.MRAM[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7907_ (.D(_0133_),
    .CLK(net235),
    .Q(\mod.Data_Mem.F_M.MRAM[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7908_ (.D(_0134_),
    .CLK(net242),
    .Q(\mod.Data_Mem.F_M.MRAM[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7909_ (.D(_0135_),
    .CLK(net236),
    .Q(\mod.Data_Mem.F_M.MRAM[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7910_ (.D(_0136_),
    .CLK(net308),
    .Q(\mod.Data_Mem.F_M.MRAM[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7911_ (.D(_0137_),
    .CLK(net368),
    .Q(\mod.Data_Mem.F_M.MRAM[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7912_ (.D(_0138_),
    .CLK(net205),
    .Q(\mod.Data_Mem.F_M.MRAM[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7913_ (.D(_0139_),
    .CLK(net155),
    .Q(\mod.Data_Mem.F_M.MRAM[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7914_ (.D(_0140_),
    .CLK(net382),
    .Q(\mod.Data_Mem.F_M.MRAM[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7915_ (.D(_0141_),
    .CLK(net368),
    .Q(\mod.Data_Mem.F_M.MRAM[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7916_ (.D(_0142_),
    .CLK(net172),
    .Q(\mod.Data_Mem.F_M.MRAM[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7917_ (.D(_0143_),
    .CLK(net174),
    .Q(\mod.Data_Mem.F_M.MRAM[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7918_ (.D(_0144_),
    .CLK(net207),
    .Q(\mod.Data_Mem.F_M.MRAM[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7919_ (.D(_0145_),
    .CLK(net201),
    .Q(\mod.Data_Mem.F_M.MRAM[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7920_ (.D(_0146_),
    .CLK(net204),
    .Q(\mod.Data_Mem.F_M.MRAM[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7921_ (.D(_0147_),
    .CLK(net209),
    .Q(\mod.Data_Mem.F_M.MRAM[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7922_ (.D(_0148_),
    .CLK(net125),
    .Q(\mod.Data_Mem.F_M.MRAM[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7923_ (.D(_0149_),
    .CLK(net122),
    .Q(\mod.Data_Mem.F_M.MRAM[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7924_ (.D(_0150_),
    .CLK(net123),
    .Q(\mod.Data_Mem.F_M.MRAM[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7925_ (.D(_0151_),
    .CLK(net125),
    .Q(\mod.Data_Mem.F_M.MRAM[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7926_ (.D(_0152_),
    .CLK(net157),
    .Q(\mod.Data_Mem.F_M.MRAM[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7927_ (.D(_0153_),
    .CLK(net372),
    .Q(\mod.Data_Mem.F_M.MRAM[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7928_ (.D(_0154_),
    .CLK(net303),
    .Q(\mod.Data_Mem.F_M.MRAM[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7929_ (.D(_0155_),
    .CLK(net368),
    .Q(\mod.Data_Mem.F_M.MRAM[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7930_ (.D(_0156_),
    .CLK(net171),
    .Q(\mod.Data_Mem.F_M.MRAM[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7931_ (.D(_0157_),
    .CLK(net386),
    .Q(\mod.Data_Mem.F_M.MRAM[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7932_ (.D(_0158_),
    .CLK(net377),
    .Q(\mod.Data_Mem.F_M.MRAM[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7933_ (.D(_0159_),
    .CLK(net166),
    .Q(\mod.Data_Mem.F_M.MRAM[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7934_ (.D(_0160_),
    .CLK(net332),
    .Q(\mod.Data_Mem.F_M.MRAM[799][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7935_ (.D(_0161_),
    .CLK(net339),
    .Q(\mod.Data_Mem.F_M.MRAM[799][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7936_ (.D(_0162_),
    .CLK(net341),
    .Q(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7937_ (.D(_0163_),
    .CLK(net288),
    .Q(\mod.Data_Mem.F_M.MRAM[799][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7938_ (.D(_0164_),
    .CLK(net97),
    .Q(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7939_ (.D(_0165_),
    .CLK(net100),
    .Q(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7940_ (.D(_0166_),
    .CLK(net98),
    .Q(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7941_ (.D(_0167_),
    .CLK(net98),
    .Q(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7942_ (.D(_0168_),
    .CLK(net138),
    .Q(\mod.Data_Mem.F_M.MRAM[789][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7943_ (.D(_0169_),
    .CLK(net154),
    .Q(\mod.Data_Mem.F_M.MRAM[789][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7944_ (.D(_0170_),
    .CLK(net190),
    .Q(\mod.Data_Mem.F_M.MRAM[789][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7945_ (.D(_0171_),
    .CLK(net142),
    .Q(\mod.Data_Mem.F_M.MRAM[789][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7946_ (.D(_0172_),
    .CLK(net88),
    .Q(\mod.Data_Mem.F_M.MRAM[789][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7947_ (.D(_0173_),
    .CLK(net138),
    .Q(\mod.Data_Mem.F_M.MRAM[789][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7948_ (.D(_0174_),
    .CLK(net85),
    .Q(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7949_ (.D(_0175_),
    .CLK(net88),
    .Q(\mod.Data_Mem.F_M.MRAM[789][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7950_ (.D(_0176_),
    .CLK(net187),
    .Q(\mod.Data_Mem.F_M.MRAM[769][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7951_ (.D(_0177_),
    .CLK(net187),
    .Q(\mod.Data_Mem.F_M.MRAM[769][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7952_ (.D(_0178_),
    .CLK(net201),
    .Q(\mod.Data_Mem.F_M.MRAM[769][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7953_ (.D(_0179_),
    .CLK(net202),
    .Q(\mod.Data_Mem.F_M.MRAM[769][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7954_ (.D(_0180_),
    .CLK(net135),
    .Q(\mod.Data_Mem.F_M.MRAM[769][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7955_ (.D(_0181_),
    .CLK(net122),
    .Q(\mod.Data_Mem.F_M.MRAM[769][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7956_ (.D(_0182_),
    .CLK(net135),
    .Q(\mod.Data_Mem.F_M.MRAM[769][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7957_ (.D(_0183_),
    .CLK(net231),
    .Q(\mod.Data_Mem.F_M.MRAM[769][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7958_ (.D(_0184_),
    .CLK(net382),
    .Q(\mod.Data_Mem.F_M.MRAM[779][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7959_ (.D(_0185_),
    .CLK(net322),
    .Q(\mod.Data_Mem.F_M.MRAM[779][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7960_ (.D(_0186_),
    .CLK(net161),
    .Q(\mod.Data_Mem.F_M.MRAM[779][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7961_ (.D(_0187_),
    .CLK(net197),
    .Q(\mod.Data_Mem.F_M.MRAM[779][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7962_ (.D(_0188_),
    .CLK(net316),
    .Q(\mod.Data_Mem.F_M.MRAM[779][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7963_ (.D(_0189_),
    .CLK(net156),
    .Q(\mod.Data_Mem.F_M.MRAM[779][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7964_ (.D(_0190_),
    .CLK(net167),
    .Q(\mod.Data_Mem.F_M.MRAM[779][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7965_ (.D(_0191_),
    .CLK(net369),
    .Q(\mod.Data_Mem.F_M.MRAM[779][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7966_ (.D(_0192_),
    .CLK(net164),
    .Q(\mod.Data_Mem.F_M.MRAM[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7967_ (.D(_0193_),
    .CLK(net144),
    .Q(\mod.Data_Mem.F_M.MRAM[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7968_ (.D(_0194_),
    .CLK(net140),
    .Q(\mod.Data_Mem.F_M.MRAM[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7969_ (.D(_0195_),
    .CLK(net163),
    .Q(\mod.Data_Mem.F_M.MRAM[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7970_ (.D(_0196_),
    .CLK(net79),
    .Q(\mod.Data_Mem.F_M.MRAM[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7971_ (.D(_0197_),
    .CLK(net158),
    .Q(\mod.Data_Mem.F_M.MRAM[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7972_ (.D(_0198_),
    .CLK(net80),
    .Q(\mod.Data_Mem.F_M.MRAM[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7973_ (.D(_0199_),
    .CLK(net72),
    .Q(\mod.Data_Mem.F_M.MRAM[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7974_ (.D(_0200_),
    .CLK(net170),
    .Q(\mod.Data_Mem.F_M.MRAM[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7975_ (.D(_0201_),
    .CLK(net149),
    .Q(\mod.Data_Mem.F_M.MRAM[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7976_ (.D(_0202_),
    .CLK(net151),
    .Q(\mod.Data_Mem.F_M.MRAM[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7977_ (.D(_0203_),
    .CLK(net184),
    .Q(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7978_ (.D(_0204_),
    .CLK(net81),
    .Q(\mod.Data_Mem.F_M.MRAM[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7979_ (.D(_0205_),
    .CLK(net89),
    .Q(\mod.Data_Mem.F_M.MRAM[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7980_ (.D(_0206_),
    .CLK(net86),
    .Q(\mod.Data_Mem.F_M.MRAM[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7981_ (.D(_0207_),
    .CLK(net81),
    .Q(\mod.Data_Mem.F_M.MRAM[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7982_ (.D(\mod.Instr_Mem.instruction[7] ),
    .RN(net25),
    .CLK(net263),
    .Q(\mod.P1.instr_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7983_ (.D(\mod.Instr_Mem.instruction[8] ),
    .RN(net34),
    .CLK(net263),
    .Q(\mod.P1.instr_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7984_ (.D(\mod.Instr_Mem.instruction[9] ),
    .RN(net16),
    .CLK(net218),
    .Q(\mod.P1.instr_reg[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7985_ (.D(\mod.Instr_Mem.instruction[10] ),
    .RN(net18),
    .CLK(net218),
    .Q(\mod.P1.instr_reg[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7986_ (.D(\mod.Instr_Mem.instruction[11] ),
    .RN(net16),
    .CLK(net219),
    .Q(\mod.P1.instr_reg[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7987_ (.D(\mod.Instr_Mem.instruction[13] ),
    .RN(net16),
    .CLK(net219),
    .Q(\mod.P1.instr_reg[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7988_ (.D(\mod.Instr_Mem.instruction[17] ),
    .RN(net21),
    .CLK(net226),
    .Q(\mod.P1.instr_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7989_ (.D(\mod.Instr_Mem.instruction[22] ),
    .RN(net11),
    .CLK(net100),
    .Q(\mod.Data_Mem.F_M.src[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7990_ (.D(\mod.Instr_Mem.instruction[23] ),
    .RN(net11),
    .CLK(net100),
    .Q(\mod.Data_Mem.F_M.src[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7991_ (.D(\mod.Instr_Mem.instruction[24] ),
    .RN(net11),
    .CLK(net115),
    .Q(\mod.Data_Mem.F_M.src[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7992_ (.D(\mod.Instr_Mem.instruction[26] ),
    .RN(net13),
    .CLK(net114),
    .Q(\mod.Data_Mem.F_M.src[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7993_ (.D(\mod.Instr_Mem.instruction[30] ),
    .RN(net18),
    .CLK(net224),
    .Q(\mod.Data_Mem.F_M.src[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7994_ (.D(\mod.P2.dest_reg1[0] ),
    .RN(net17),
    .CLK(net223),
    .Q(\mod.P2.dest_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7995_ (.D(\mod.P2.dest_reg1[1] ),
    .RN(net19),
    .CLK(net226),
    .Q(\mod.P2.dest_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7996_ (.D(\mod.P2.dest_reg1[2] ),
    .RN(net20),
    .CLK(net224),
    .Q(\mod.P2.dest_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7997_ (.D(\mod.P2.dest_reg1[4] ),
    .RN(net20),
    .CLK(net223),
    .Q(\mod.P2.dest_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _7998_ (.D(\mod.P2.dest_reg1[8] ),
    .RN(net25),
    .CLK(net240),
    .Q(\mod.P2.dest_reg[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7999_ (.D(_0208_),
    .CLK(net305),
    .Q(\mod.Data_Mem.F_M.MRAM[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8000_ (.D(_0209_),
    .CLK(net297),
    .Q(\mod.Data_Mem.F_M.MRAM[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8001_ (.D(_0210_),
    .CLK(net297),
    .Q(\mod.Data_Mem.F_M.MRAM[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8002_ (.D(_0211_),
    .CLK(net305),
    .Q(\mod.Data_Mem.F_M.MRAM[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8003_ (.D(_0212_),
    .CLK(net232),
    .Q(\mod.Data_Mem.F_M.MRAM[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8004_ (.D(_0213_),
    .CLK(net232),
    .Q(\mod.Data_Mem.F_M.MRAM[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8005_ (.D(_0214_),
    .CLK(net259),
    .Q(\mod.Data_Mem.F_M.MRAM[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8006_ (.D(_0215_),
    .CLK(net233),
    .Q(\mod.Data_Mem.F_M.MRAM[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8007_ (.D(_0216_),
    .CLK(net301),
    .Q(\mod.Data_Mem.F_M.MRAM[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8008_ (.D(_0217_),
    .CLK(net302),
    .Q(\mod.Data_Mem.F_M.MRAM[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8009_ (.D(_0218_),
    .CLK(net305),
    .Q(\mod.Data_Mem.F_M.MRAM[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8010_ (.D(_0219_),
    .CLK(net305),
    .Q(\mod.Data_Mem.F_M.MRAM[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8011_ (.D(_0220_),
    .CLK(net233),
    .Q(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8012_ (.D(_0221_),
    .CLK(net231),
    .Q(\mod.Data_Mem.F_M.MRAM[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8013_ (.D(_0222_),
    .CLK(net126),
    .Q(\mod.Data_Mem.F_M.MRAM[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8014_ (.D(_0223_),
    .CLK(net126),
    .Q(\mod.Data_Mem.F_M.MRAM[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8015_ (.D(_0224_),
    .CLK(net303),
    .Q(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8016_ (.D(_0225_),
    .CLK(net302),
    .Q(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8017_ (.D(_0226_),
    .CLK(net306),
    .Q(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8018_ (.D(_0227_),
    .CLK(net306),
    .Q(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8019_ (.D(_0228_),
    .CLK(net232),
    .Q(\mod.Data_Mem.F_M.MRAM[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8020_ (.D(_0229_),
    .CLK(net109),
    .Q(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8021_ (.D(_0230_),
    .CLK(net109),
    .Q(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8022_ (.D(_0231_),
    .CLK(net122),
    .Q(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8023_ (.D(_0232_),
    .CLK(net210),
    .Q(\mod.Data_Mem.F_M.MRAM[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8024_ (.D(_0233_),
    .CLK(net301),
    .Q(\mod.Data_Mem.F_M.MRAM[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8025_ (.D(_0234_),
    .CLK(net301),
    .Q(\mod.Data_Mem.F_M.MRAM[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8026_ (.D(_0235_),
    .CLK(net209),
    .Q(\mod.Data_Mem.F_M.MRAM[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8027_ (.D(_0236_),
    .CLK(net70),
    .Q(\mod.Data_Mem.F_M.MRAM[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8028_ (.D(_0237_),
    .CLK(net70),
    .Q(\mod.Data_Mem.F_M.MRAM[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8029_ (.D(_0238_),
    .CLK(net73),
    .Q(\mod.Data_Mem.F_M.MRAM[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8030_ (.D(_0239_),
    .CLK(net73),
    .Q(\mod.Data_Mem.F_M.MRAM[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8031_ (.D(_0240_),
    .CLK(net210),
    .Q(\mod.Data_Mem.F_M.MRAM[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8032_ (.D(_0241_),
    .CLK(net211),
    .Q(\mod.Data_Mem.F_M.MRAM[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8033_ (.D(_0242_),
    .CLK(net301),
    .Q(\mod.Data_Mem.F_M.MRAM[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8034_ (.D(_0243_),
    .CLK(net210),
    .Q(\mod.Data_Mem.F_M.MRAM[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8035_ (.D(_0244_),
    .CLK(net71),
    .Q(\mod.Data_Mem.F_M.MRAM[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8036_ (.D(_0245_),
    .CLK(net70),
    .Q(\mod.Data_Mem.F_M.MRAM[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8037_ (.D(_0246_),
    .CLK(net73),
    .Q(\mod.Data_Mem.F_M.MRAM[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8038_ (.D(_0247_),
    .CLK(net74),
    .Q(\mod.Data_Mem.F_M.MRAM[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8039_ (.D(_0248_),
    .CLK(net191),
    .Q(\mod.Data_Mem.F_M.MRAM[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8040_ (.D(_0249_),
    .CLK(net195),
    .Q(\mod.Data_Mem.F_M.MRAM[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8041_ (.D(_0250_),
    .CLK(net195),
    .Q(\mod.Data_Mem.F_M.MRAM[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8042_ (.D(_0251_),
    .CLK(net195),
    .Q(\mod.Data_Mem.F_M.MRAM[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8043_ (.D(_0252_),
    .CLK(net71),
    .Q(\mod.Data_Mem.F_M.MRAM[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8044_ (.D(_0253_),
    .CLK(net78),
    .Q(\mod.Data_Mem.F_M.MRAM[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8045_ (.D(_0254_),
    .CLK(net106),
    .Q(\mod.Data_Mem.F_M.MRAM[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8046_ (.D(_0255_),
    .CLK(net106),
    .Q(\mod.Data_Mem.F_M.MRAM[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8047_ (.D(_0256_),
    .CLK(net207),
    .Q(\mod.Data_Mem.F_M.MRAM[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8048_ (.D(_0257_),
    .CLK(net207),
    .Q(\mod.Data_Mem.F_M.MRAM[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8049_ (.D(_0258_),
    .CLK(net209),
    .Q(\mod.Data_Mem.F_M.MRAM[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8050_ (.D(_0259_),
    .CLK(net209),
    .Q(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8051_ (.D(_0260_),
    .CLK(net125),
    .Q(\mod.Data_Mem.F_M.MRAM[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8052_ (.D(_0261_),
    .CLK(net123),
    .Q(\mod.Data_Mem.F_M.MRAM[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8053_ (.D(_0262_),
    .CLK(net123),
    .Q(\mod.Data_Mem.F_M.MRAM[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8054_ (.D(_0263_),
    .CLK(net125),
    .Q(\mod.Data_Mem.F_M.MRAM[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8055_ (.D(_0264_),
    .CLK(net163),
    .Q(\mod.Data_Mem.F_M.MRAM[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8056_ (.D(_0265_),
    .CLK(net147),
    .Q(\mod.Data_Mem.F_M.MRAM[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8057_ (.D(_0266_),
    .CLK(net147),
    .Q(\mod.Data_Mem.F_M.MRAM[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8058_ (.D(_0267_),
    .CLK(net184),
    .Q(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8059_ (.D(_0268_),
    .CLK(net95),
    .Q(\mod.Data_Mem.F_M.MRAM[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8060_ (.D(_0269_),
    .CLK(net89),
    .Q(\mod.Data_Mem.F_M.MRAM[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8061_ (.D(_0270_),
    .CLK(net75),
    .Q(\mod.Data_Mem.F_M.MRAM[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8062_ (.D(_0271_),
    .CLK(net80),
    .Q(\mod.Data_Mem.F_M.MRAM[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8063_ (.D(_0272_),
    .CLK(net163),
    .Q(\mod.Data_Mem.F_M.MRAM[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8064_ (.D(_0273_),
    .CLK(net147),
    .Q(\mod.Data_Mem.F_M.MRAM[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8065_ (.D(_0274_),
    .CLK(net148),
    .Q(\mod.Data_Mem.F_M.MRAM[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8066_ (.D(_0275_),
    .CLK(net186),
    .Q(\mod.Data_Mem.F_M.MRAM[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8067_ (.D(_0276_),
    .CLK(net82),
    .Q(\mod.Data_Mem.F_M.MRAM[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8068_ (.D(_0277_),
    .CLK(net91),
    .Q(\mod.Data_Mem.F_M.MRAM[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8069_ (.D(_0278_),
    .CLK(net75),
    .Q(\mod.Data_Mem.F_M.MRAM[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8070_ (.D(_0279_),
    .CLK(net132),
    .Q(\mod.Data_Mem.F_M.MRAM[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8071_ (.D(\mod.DMen_reg ),
    .RN(net25),
    .CLK(net237),
    .Q(\mod.DMen_reg2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8072_ (.D(\mod.P3.Res[0] ),
    .RN(net61),
    .CLK(net384),
    .Q(net3));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8073_ (.D(\mod.P3.Res[1] ),
    .RN(net32),
    .CLK(net246),
    .Q(net4));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8074_ (.D(\mod.P3.Res[2] ),
    .RN(net36),
    .CLK(net284),
    .Q(net5));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8075_ (.D(\mod.P3.Res[3] ),
    .RN(net32),
    .CLK(net245),
    .Q(net6));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8076_ (.D(\mod.P3.Res[4] ),
    .RN(net34),
    .CLK(net261),
    .Q(net7));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8077_ (.D(\mod.P3.Res[5] ),
    .RN(net26),
    .CLK(net264),
    .Q(net8));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8078_ (.D(\mod.P3.Res[6] ),
    .RN(net34),
    .CLK(net262),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8079_ (.D(\mod.P3.Res[7] ),
    .RN(net26),
    .CLK(net245),
    .Q(net10));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8080_ (.D(_0280_),
    .CLK(net160),
    .Q(\mod.Data_Mem.F_M.MRAM[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8081_ (.D(_0281_),
    .CLK(net140),
    .Q(\mod.Data_Mem.F_M.MRAM[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8082_ (.D(_0282_),
    .CLK(net141),
    .Q(\mod.Data_Mem.F_M.MRAM[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8083_ (.D(_0283_),
    .CLK(net304),
    .Q(\mod.Data_Mem.F_M.MRAM[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8084_ (.D(_0284_),
    .CLK(net73),
    .Q(\mod.Data_Mem.F_M.MRAM[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8085_ (.D(_0285_),
    .CLK(net88),
    .Q(\mod.Data_Mem.F_M.MRAM[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8086_ (.D(_0286_),
    .CLK(net78),
    .Q(\mod.Data_Mem.F_M.MRAM[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8087_ (.D(_0287_),
    .CLK(net81),
    .Q(\mod.Data_Mem.F_M.MRAM[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8088_ (.D(\mod.P2.Rout_reg1[0] ),
    .RN(net35),
    .CLK(net261),
    .Q(\mod.P2.Rout_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8089_ (.D(\mod.P2.Rout_reg1[1] ),
    .RN(net35),
    .CLK(net261),
    .Q(\mod.P2.Rout_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8090_ (.D(\mod.Data_Mem.F_M.out_data[0] ),
    .RN(net54),
    .CLK(net344),
    .Q(\mod.Arithmetic.ACTI.x[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8091_ (.D(\mod.Data_Mem.F_M.out_data[1] ),
    .RN(net58),
    .CLK(net345),
    .Q(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8092_ (.D(\mod.Data_Mem.F_M.out_data[2] ),
    .RN(net59),
    .CLK(net348),
    .Q(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8093_ (.D(\mod.Data_Mem.F_M.out_data[3] ),
    .RN(net56),
    .CLK(net336),
    .Q(\mod.Arithmetic.ACTI.x[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8094_ (.D(\mod.Data_Mem.F_M.out_data[4] ),
    .RN(net28),
    .CLK(net268),
    .Q(\mod.Arithmetic.ACTI.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8095_ (.D(\mod.Data_Mem.F_M.out_data[5] ),
    .RN(net51),
    .CLK(net282),
    .Q(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8096_ (.D(\mod.Data_Mem.F_M.out_data[6] ),
    .RN(net26),
    .CLK(net266),
    .Q(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8097_ (.D(\mod.Data_Mem.F_M.out_data[7] ),
    .RN(net26),
    .CLK(net246),
    .Q(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8098_ (.D(\mod.Data_Mem.F_M.out_data[8] ),
    .RN(net55),
    .CLK(net345),
    .Q(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8099_ (.D(\mod.Data_Mem.F_M.out_data[9] ),
    .RN(net52),
    .CLK(net344),
    .Q(\mod.Arithmetic.CN.I_in[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8100_ (.D(\mod.Data_Mem.F_M.out_data[10] ),
    .RN(net58),
    .CLK(net345),
    .Q(\mod.Arithmetic.CN.I_in[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8101_ (.D(\mod.Data_Mem.F_M.out_data[11] ),
    .RN(net36),
    .CLK(net282),
    .Q(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8102_ (.D(\mod.Data_Mem.F_M.out_data[12] ),
    .RN(net32),
    .CLK(net247),
    .Q(\mod.Arithmetic.CN.I_in[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8103_ (.D(\mod.Data_Mem.F_M.out_data[13] ),
    .RN(net30),
    .CLK(net270),
    .Q(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8104_ (.D(\mod.Data_Mem.F_M.out_data[14] ),
    .RN(net30),
    .CLK(net269),
    .Q(\mod.Arithmetic.CN.I_in[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8105_ (.D(\mod.Data_Mem.F_M.out_data[15] ),
    .RN(net28),
    .CLK(net268),
    .Q(\mod.Arithmetic.CN.I_in[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8106_ (.D(\mod.Data_Mem.F_M.out_data[16] ),
    .RN(net42),
    .CLK(net275),
    .Q(\mod.Arithmetic.CN.I_in[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8107_ (.D(\mod.Data_Mem.F_M.out_data[17] ),
    .RN(net54),
    .CLK(net341),
    .Q(\mod.Arithmetic.CN.I_in[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8108_ (.D(\mod.Data_Mem.F_M.out_data[18] ),
    .RN(net54),
    .CLK(net349),
    .Q(\mod.Arithmetic.CN.I_in[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8109_ (.D(\mod.Data_Mem.F_M.out_data[19] ),
    .RN(net46),
    .CLK(net329),
    .Q(\mod.Arithmetic.CN.I_in[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8110_ (.D(\mod.Data_Mem.F_M.out_data[20] ),
    .RN(net42),
    .CLK(net278),
    .Q(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8111_ (.D(\mod.Data_Mem.F_M.out_data[21] ),
    .RN(net43),
    .CLK(net278),
    .Q(\mod.Arithmetic.CN.I_in[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8112_ (.D(\mod.Data_Mem.F_M.out_data[22] ),
    .RN(net40),
    .CLK(net274),
    .Q(\mod.Arithmetic.CN.I_in[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8113_ (.D(\mod.Data_Mem.F_M.out_data[23] ),
    .RN(net40),
    .CLK(net274),
    .Q(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8114_ (.D(\mod.Data_Mem.F_M.out_data[24] ),
    .RN(net46),
    .CLK(net329),
    .Q(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8115_ (.D(\mod.Data_Mem.F_M.out_data[25] ),
    .RN(net51),
    .CLK(net337),
    .Q(\mod.Arithmetic.CN.I_in[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8116_ (.D(\mod.Data_Mem.F_M.out_data[26] ),
    .RN(net52),
    .CLK(net334),
    .Q(\mod.Arithmetic.CN.I_in[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8117_ (.D(\mod.Data_Mem.F_M.out_data[27] ),
    .RN(net46),
    .CLK(net329),
    .Q(\mod.Arithmetic.CN.I_in[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8118_ (.D(\mod.Data_Mem.F_M.out_data[28] ),
    .RN(net41),
    .CLK(net274),
    .Q(\mod.Arithmetic.CN.I_in[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8119_ (.D(\mod.Data_Mem.F_M.out_data[29] ),
    .RN(net43),
    .CLK(net278),
    .Q(\mod.Arithmetic.CN.I_in[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8120_ (.D(\mod.Data_Mem.F_M.out_data[30] ),
    .RN(net41),
    .CLK(net276),
    .Q(\mod.Arithmetic.CN.I_in[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8121_ (.D(\mod.Data_Mem.F_M.out_data[31] ),
    .RN(net40),
    .CLK(net274),
    .Q(\mod.Arithmetic.CN.I_in[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8122_ (.D(\mod.Data_Mem.F_M.out_data[32] ),
    .RN(net48),
    .CLK(net337),
    .Q(\mod.Arithmetic.CN.I_in[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8123_ (.D(\mod.Data_Mem.F_M.out_data[33] ),
    .RN(net58),
    .CLK(net346),
    .Q(\mod.Arithmetic.CN.I_in[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8124_ (.D(\mod.Data_Mem.F_M.out_data[34] ),
    .RN(net59),
    .CLK(net355),
    .Q(\mod.Arithmetic.CN.I_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8125_ (.D(\mod.Data_Mem.F_M.out_data[35] ),
    .RN(net47),
    .CLK(net278),
    .Q(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8126_ (.D(\mod.Data_Mem.F_M.out_data[36] ),
    .RN(net30),
    .CLK(net273),
    .Q(\mod.Arithmetic.CN.I_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8127_ (.D(\mod.Data_Mem.F_M.out_data[37] ),
    .RN(net37),
    .CLK(net273),
    .Q(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8128_ (.D(\mod.Data_Mem.F_M.out_data[38] ),
    .RN(net44),
    .CLK(net251),
    .Q(\mod.Arithmetic.CN.I_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8129_ (.D(\mod.Data_Mem.F_M.out_data[39] ),
    .RN(net40),
    .CLK(net275),
    .Q(\mod.Arithmetic.CN.I_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8130_ (.D(\mod.Data_Mem.F_M.out_data[40] ),
    .RN(net51),
    .CLK(net334),
    .Q(\mod.Arithmetic.CN.I_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8131_ (.D(\mod.Data_Mem.F_M.out_data[41] ),
    .RN(net52),
    .CLK(net330),
    .Q(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8132_ (.D(\mod.Data_Mem.F_M.out_data[42] ),
    .RN(net46),
    .CLK(net327),
    .Q(\mod.Arithmetic.CN.I_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8133_ (.D(\mod.Data_Mem.F_M.out_data[43] ),
    .RN(net47),
    .CLK(net279),
    .Q(\mod.Arithmetic.CN.I_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8134_ (.D(\mod.Data_Mem.F_M.out_data[44] ),
    .RN(net44),
    .CLK(net255),
    .Q(\mod.Arithmetic.CN.I_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8135_ (.D(\mod.Data_Mem.F_M.out_data[45] ),
    .RN(net47),
    .CLK(net279),
    .Q(\mod.Arithmetic.CN.I_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8136_ (.D(\mod.Data_Mem.F_M.out_data[46] ),
    .RN(net44),
    .CLK(net251),
    .Q(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8137_ (.D(\mod.Data_Mem.F_M.out_data[47] ),
    .RN(net44),
    .CLK(net255),
    .Q(\mod.Arithmetic.CN.I_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8138_ (.D(\mod.Data_Mem.F_M.out_data[48] ),
    .RN(net59),
    .CLK(net348),
    .Q(\mod.Arithmetic.CN.I_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8139_ (.D(\mod.Data_Mem.F_M.out_data[49] ),
    .RN(net53),
    .CLK(net331),
    .Q(\mod.Arithmetic.CN.I_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8140_ (.D(\mod.Data_Mem.F_M.out_data[50] ),
    .RN(net55),
    .CLK(net354),
    .Q(\mod.Arithmetic.CN.I_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8141_ (.D(\mod.Data_Mem.F_M.out_data[51] ),
    .RN(net55),
    .CLK(net354),
    .Q(\mod.Arithmetic.CN.I_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8142_ (.D(\mod.Data_Mem.F_M.out_data[52] ),
    .RN(net63),
    .CLK(net354),
    .Q(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8143_ (.D(\mod.Data_Mem.F_M.out_data[53] ),
    .RN(net63),
    .CLK(net356),
    .Q(\mod.Arithmetic.CN.I_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8144_ (.D(\mod.Data_Mem.F_M.out_data[54] ),
    .RN(net63),
    .CLK(net363),
    .Q(\mod.Arithmetic.CN.I_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8145_ (.D(\mod.Data_Mem.F_M.out_data[55] ),
    .RN(net63),
    .CLK(net361),
    .Q(\mod.Arithmetic.CN.I_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8146_ (.D(\mod.Data_Mem.F_M.out_data[56] ),
    .RN(net67),
    .CLK(net344),
    .Q(\mod.Arithmetic.CN.I_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8147_ (.D(\mod.Data_Mem.F_M.out_data[57] ),
    .RN(net52),
    .CLK(net334),
    .Q(\mod.Arithmetic.CN.I_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8148_ (.D(\mod.Data_Mem.F_M.out_data[58] ),
    .RN(net55),
    .CLK(net335),
    .Q(\mod.Arithmetic.CN.I_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8149_ (.D(\mod.Data_Mem.F_M.out_data[59] ),
    .RN(net57),
    .CLK(net354),
    .Q(\mod.Arithmetic.CN.I_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8150_ (.D(\mod.Data_Mem.F_M.out_data[60] ),
    .RN(net62),
    .CLK(net363),
    .Q(\mod.Arithmetic.CN.I_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8151_ (.D(\mod.Data_Mem.F_M.out_data[61] ),
    .RN(net61),
    .CLK(net361),
    .Q(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8152_ (.D(\mod.Data_Mem.F_M.out_data[62] ),
    .RN(net61),
    .CLK(net362),
    .Q(\mod.Arithmetic.CN.I_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8153_ (.D(\mod.Data_Mem.F_M.out_data[63] ),
    .RN(net61),
    .CLK(net361),
    .Q(\mod.Arithmetic.CN.I_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8154_ (.D(\mod.Data_Mem.F_M.out_data[64] ),
    .RN(net60),
    .CLK(net348),
    .Q(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8155_ (.D(\mod.Data_Mem.F_M.out_data[65] ),
    .RN(net56),
    .CLK(net336),
    .Q(\mod.Arithmetic.CN.I_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8156_ (.D(\mod.Data_Mem.F_M.out_data[66] ),
    .RN(net58),
    .CLK(net357),
    .Q(\mod.Arithmetic.CN.I_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8157_ (.D(\mod.Data_Mem.F_M.out_data[67] ),
    .RN(net56),
    .CLK(net355),
    .Q(\mod.Arithmetic.CN.I_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8158_ (.D(\mod.Data_Mem.F_M.out_data[68] ),
    .RN(net60),
    .CLK(net358),
    .Q(\mod.Arithmetic.CN.I_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8159_ (.D(\mod.Data_Mem.F_M.out_data[69] ),
    .RN(net62),
    .CLK(net358),
    .Q(\mod.Arithmetic.CN.I_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8160_ (.D(\mod.Data_Mem.F_M.out_data[70] ),
    .RN(net64),
    .CLK(net383),
    .Q(\mod.Arithmetic.CN.I_in[70] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8161_ (.D(\mod.Data_Mem.F_M.out_data[71] ),
    .RN(net62),
    .CLK(net358),
    .Q(\mod.Arithmetic.CN.I_in[71] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8162_ (.D(\mod.Data_Mem.F_M.out_data[72] ),
    .RN(net30),
    .CLK(net270),
    .Q(\mod.Arithmetic.I_out[72] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8163_ (.D(\mod.Data_Mem.F_M.out_data[73] ),
    .RN(net29),
    .CLK(net270),
    .Q(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8164_ (.D(\mod.Data_Mem.F_M.out_data[74] ),
    .RN(net31),
    .CLK(net270),
    .Q(\mod.Arithmetic.I_out[74] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8165_ (.D(\mod.Data_Mem.F_M.out_data[75] ),
    .RN(net28),
    .CLK(net266),
    .Q(\mod.Arithmetic.I_out[75] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8166_ (.D(\mod.Data_Mem.F_M.out_data[76] ),
    .RN(net28),
    .CLK(net266),
    .Q(\mod.Arithmetic.I_out[76] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8167_ (.D(\mod.Data_Mem.F_M.out_data[77] ),
    .RN(net29),
    .CLK(net267),
    .Q(\mod.Arithmetic.I_out[77] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _8168_ (.D(\mod.Data_Mem.F_M.out_data[78] ),
    .RN(net27),
    .CLK(net266),
    .Q(\mod.Arithmetic.I_out[78] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8169_ (.D(\mod.Data_Mem.F_M.out_data[79] ),
    .RN(net27),
    .CLK(net264),
    .Q(\mod.Arithmetic.I_out[79] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8170_ (.D(\mod.P2.dest_reg[0] ),
    .RN(net20),
    .CLK(net223),
    .Q(\mod.Data_Mem.F_M.dest[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8171_ (.D(\mod.P2.dest_reg[1] ),
    .RN(net21),
    .CLK(net227),
    .Q(\mod.Data_Mem.F_M.dest[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8172_ (.D(\mod.P2.dest_reg[2] ),
    .RN(net21),
    .CLK(net225),
    .Q(\mod.Data_Mem.F_M.dest[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8173_ (.D(\mod.P2.dest_reg[4] ),
    .RN(net20),
    .CLK(net225),
    .Q(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8174_ (.D(\mod.P2.dest_reg[8] ),
    .RN(net25),
    .CLK(net237),
    .Q(\mod.Data_Mem.F_M.dest[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8175_ (.D(\mod.DM_en ),
    .RN(net23),
    .CLK(net235),
    .Q(\mod.DMen_reg ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8176_ (.D(\mod.P1.instr_reg[7] ),
    .RN(net38),
    .CLK(net262),
    .Q(\mod.P2.Rout_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8177_ (.D(\mod.P1.instr_reg[8] ),
    .RN(net34),
    .CLK(net261),
    .Q(\mod.P2.Rout_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8178_ (.D(_0288_),
    .CLK(net191),
    .Q(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8179_ (.D(_0289_),
    .CLK(net206),
    .Q(\mod.Data_Mem.F_M.MRAM[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8180_ (.D(_0290_),
    .CLK(net207),
    .Q(\mod.Data_Mem.F_M.MRAM[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8181_ (.D(_0291_),
    .CLK(net206),
    .Q(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8182_ (.D(_0292_),
    .CLK(net109),
    .Q(\mod.Data_Mem.F_M.MRAM[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8183_ (.D(_0293_),
    .CLK(net106),
    .Q(\mod.Data_Mem.F_M.MRAM[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8184_ (.D(_0294_),
    .CLK(net76),
    .Q(\mod.Data_Mem.F_M.MRAM[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8185_ (.D(_0295_),
    .CLK(net107),
    .Q(\mod.Data_Mem.F_M.MRAM[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8186_ (.D(_0296_),
    .CLK(net191),
    .Q(\mod.Data_Mem.F_M.MRAM[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8187_ (.D(_0297_),
    .CLK(net196),
    .Q(\mod.Data_Mem.F_M.MRAM[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8188_ (.D(_0298_),
    .CLK(net195),
    .Q(\mod.Data_Mem.F_M.MRAM[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8189_ (.D(_0299_),
    .CLK(net196),
    .Q(\mod.Data_Mem.F_M.MRAM[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8190_ (.D(_0300_),
    .CLK(net70),
    .Q(\mod.Data_Mem.F_M.MRAM[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8191_ (.D(_0301_),
    .CLK(net78),
    .Q(\mod.Data_Mem.F_M.MRAM[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8192_ (.D(_0302_),
    .CLK(net106),
    .Q(\mod.Data_Mem.F_M.MRAM[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8193_ (.D(_0303_),
    .CLK(net109),
    .Q(\mod.Data_Mem.F_M.MRAM[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8194_ (.D(net574),
    .RN(net47),
    .CLK(net333),
    .Q(\mod.Arithmetic.CN.F_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8195_ (.D(_0080_),
    .RN(net14),
    .CLK(net118),
    .Q(\mod.I_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8196_ (.D(_0081_),
    .RN(net14),
    .CLK(net118),
    .Q(\mod.I_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8197_ (.D(_0082_),
    .RN(net15),
    .CLK(net118),
    .Q(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8198_ (.D(_0083_),
    .RN(net14),
    .CLK(net118),
    .Q(\mod.I_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8199_ (.D(_0084_),
    .RN(net14),
    .CLK(net114),
    .Q(\mod.I_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8200_ (.D(_0085_),
    .RN(net11),
    .CLK(net114),
    .Q(\mod.I_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8201_ (.D(_0086_),
    .RN(net12),
    .CLK(net114),
    .Q(\mod.I_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8202_ (.D(_0087_),
    .RN(net12),
    .CLK(net115),
    .Q(\mod.I_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8203_ (.D(_0304_),
    .CLK(net297),
    .Q(\mod.Data_Mem.F_M.MRAM[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8204_ (.D(_0305_),
    .CLK(net296),
    .Q(\mod.Data_Mem.F_M.MRAM[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8205_ (.D(_0306_),
    .CLK(net297),
    .Q(\mod.Data_Mem.F_M.MRAM[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8206_ (.D(_0307_),
    .CLK(net299),
    .Q(\mod.Data_Mem.F_M.MRAM[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8207_ (.D(_0308_),
    .CLK(net243),
    .Q(\mod.Data_Mem.F_M.MRAM[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8208_ (.D(_0309_),
    .CLK(net245),
    .Q(\mod.Data_Mem.F_M.MRAM[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8209_ (.D(_0310_),
    .CLK(net242),
    .Q(\mod.Data_Mem.F_M.MRAM[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8210_ (.D(_0311_),
    .CLK(net243),
    .Q(\mod.Data_Mem.F_M.MRAM[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8211_ (.D(_0312_),
    .CLK(net161),
    .Q(\mod.Data_Mem.F_M.MRAM[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8212_ (.D(_0313_),
    .CLK(net144),
    .Q(\mod.Data_Mem.F_M.MRAM[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8213_ (.D(_0314_),
    .CLK(net145),
    .Q(\mod.Data_Mem.F_M.MRAM[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8214_ (.D(_0315_),
    .CLK(net150),
    .Q(\mod.Data_Mem.F_M.MRAM[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8215_ (.D(_0316_),
    .CLK(net72),
    .Q(\mod.Data_Mem.F_M.MRAM[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8216_ (.D(_0317_),
    .CLK(net89),
    .Q(\mod.Data_Mem.F_M.MRAM[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8217_ (.D(_0318_),
    .CLK(net78),
    .Q(\mod.Data_Mem.F_M.MRAM[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8218_ (.D(_0319_),
    .CLK(net81),
    .Q(\mod.Data_Mem.F_M.MRAM[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8219_ (.D(_0320_),
    .CLK(net299),
    .Q(\mod.Data_Mem.F_M.MRAM[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8220_ (.D(_0321_),
    .CLK(net311),
    .Q(\mod.Data_Mem.F_M.MRAM[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8221_ (.D(_0322_),
    .CLK(net311),
    .Q(\mod.Data_Mem.F_M.MRAM[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8222_ (.D(_0323_),
    .CLK(net311),
    .Q(\mod.Data_Mem.F_M.MRAM[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8223_ (.D(_0324_),
    .CLK(net244),
    .Q(\mod.Data_Mem.F_M.MRAM[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8224_ (.D(_0325_),
    .CLK(net248),
    .Q(\mod.Data_Mem.F_M.MRAM[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8225_ (.D(_0326_),
    .CLK(net244),
    .Q(\mod.Data_Mem.F_M.MRAM[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8226_ (.D(_0327_),
    .CLK(net242),
    .Q(\mod.Data_Mem.F_M.MRAM[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8227_ (.D(\mod.P1.instr_reg[9] ),
    .RN(net16),
    .CLK(net219),
    .Q(\mod.P2.dest_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8228_ (.D(\mod.P1.instr_reg[10] ),
    .RN(net19),
    .CLK(net219),
    .Q(\mod.P2.dest_reg1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8229_ (.D(\mod.P1.instr_reg[11] ),
    .RN(net17),
    .CLK(net224),
    .Q(\mod.P2.dest_reg1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8230_ (.D(\mod.P1.instr_reg[13] ),
    .RN(net17),
    .CLK(net223),
    .Q(\mod.P2.dest_reg1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _8231_ (.D(\mod.P1.instr_reg[17] ),
    .RN(net23),
    .CLK(net240),
    .Q(\mod.P2.dest_reg1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8232_ (.D(_0328_),
    .CLK(net296),
    .Q(\mod.Data_Mem.F_M.MRAM[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8233_ (.D(_0329_),
    .CLK(net204),
    .Q(\mod.Data_Mem.F_M.MRAM[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8234_ (.D(_0330_),
    .CLK(net300),
    .Q(\mod.Data_Mem.F_M.MRAM[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8235_ (.D(_0331_),
    .CLK(net213),
    .Q(\mod.Data_Mem.F_M.MRAM[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8236_ (.D(_0332_),
    .CLK(net135),
    .Q(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8237_ (.D(_0333_),
    .CLK(net132),
    .Q(\mod.Data_Mem.F_M.MRAM[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8238_ (.D(_0334_),
    .CLK(net107),
    .Q(\mod.Data_Mem.F_M.MRAM[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8239_ (.D(_0335_),
    .CLK(net132),
    .Q(\mod.Data_Mem.F_M.MRAM[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8240_ (.D(_0336_),
    .CLK(net298),
    .Q(\mod.Data_Mem.F_M.MRAM[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8241_ (.D(_0337_),
    .CLK(net312),
    .Q(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8242_ (.D(_0338_),
    .CLK(net313),
    .Q(\mod.Data_Mem.F_M.MRAM[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8243_ (.D(_0339_),
    .CLK(net298),
    .Q(\mod.Data_Mem.F_M.MRAM[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8244_ (.D(_0340_),
    .CLK(net136),
    .Q(\mod.Data_Mem.F_M.MRAM[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8245_ (.D(_0341_),
    .CLK(net132),
    .Q(\mod.Data_Mem.F_M.MRAM[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8246_ (.D(_0342_),
    .CLK(net133),
    .Q(\mod.Data_Mem.F_M.MRAM[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8247_ (.D(_0343_),
    .CLK(net133),
    .Q(\mod.Data_Mem.F_M.MRAM[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8248_ (.D(_0344_),
    .CLK(net339),
    .Q(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8249_ (.D(_0345_),
    .CLK(net314),
    .Q(\mod.Data_Mem.F_M.MRAM[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8250_ (.D(_0346_),
    .CLK(net341),
    .Q(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8251_ (.D(_0347_),
    .CLK(net311),
    .Q(\mod.Data_Mem.F_M.MRAM[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8252_ (.D(_0348_),
    .CLK(net101),
    .Q(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8253_ (.D(_0349_),
    .CLK(net116),
    .Q(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8254_ (.D(_0350_),
    .CLK(net116),
    .Q(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8255_ (.D(_0351_),
    .CLK(net116),
    .Q(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8256_ (.D(_0352_),
    .CLK(net163),
    .Q(\mod.Data_Mem.F_M.MRAM[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8257_ (.D(_0353_),
    .CLK(net149),
    .Q(\mod.Data_Mem.F_M.MRAM[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8258_ (.D(_0354_),
    .CLK(net149),
    .Q(\mod.Data_Mem.F_M.MRAM[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8259_ (.D(_0355_),
    .CLK(net184),
    .Q(\mod.Data_Mem.F_M.MRAM[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8260_ (.D(_0356_),
    .CLK(net82),
    .Q(\mod.Data_Mem.F_M.MRAM[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8261_ (.D(_0357_),
    .CLK(net92),
    .Q(\mod.Data_Mem.F_M.MRAM[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8262_ (.D(_0358_),
    .CLK(net91),
    .Q(\mod.Data_Mem.F_M.MRAM[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8263_ (.D(_0359_),
    .CLK(net82),
    .Q(\mod.Data_Mem.F_M.MRAM[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8264_ (.D(_0360_),
    .CLK(net187),
    .Q(\mod.Data_Mem.F_M.MRAM[768][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8265_ (.D(_0361_),
    .CLK(net203),
    .Q(\mod.Data_Mem.F_M.MRAM[768][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8266_ (.D(_0362_),
    .CLK(net203),
    .Q(\mod.Data_Mem.F_M.MRAM[768][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8267_ (.D(_0363_),
    .CLK(net183),
    .Q(\mod.Data_Mem.F_M.MRAM[768][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8268_ (.D(_0364_),
    .CLK(net127),
    .Q(\mod.Data_Mem.F_M.MRAM[768][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8269_ (.D(_0365_),
    .CLK(net122),
    .Q(\mod.Data_Mem.F_M.MRAM[768][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8270_ (.D(_0366_),
    .CLK(net127),
    .Q(\mod.Data_Mem.F_M.MRAM[768][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8271_ (.D(_0367_),
    .CLK(net127),
    .Q(\mod.Data_Mem.F_M.MRAM[768][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8272_ (.D(_0368_),
    .CLK(net187),
    .Q(\mod.Data_Mem.F_M.MRAM[770][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8273_ (.D(_0369_),
    .CLK(net203),
    .Q(\mod.Data_Mem.F_M.MRAM[770][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8274_ (.D(_0370_),
    .CLK(net203),
    .Q(\mod.Data_Mem.F_M.MRAM[770][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8275_ (.D(_0371_),
    .CLK(net183),
    .Q(\mod.Data_Mem.F_M.MRAM[770][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8276_ (.D(_0372_),
    .CLK(net110),
    .Q(\mod.Data_Mem.F_M.MRAM[770][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8277_ (.D(_0373_),
    .CLK(net111),
    .Q(\mod.Data_Mem.F_M.MRAM[770][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8278_ (.D(_0374_),
    .CLK(net121),
    .Q(\mod.Data_Mem.F_M.MRAM[770][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8279_ (.D(_0375_),
    .CLK(net121),
    .Q(\mod.Data_Mem.F_M.MRAM[770][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8280_ (.D(_0376_),
    .CLK(net296),
    .Q(\mod.Data_Mem.F_M.MRAM[771][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8281_ (.D(_0377_),
    .CLK(net314),
    .Q(\mod.Data_Mem.F_M.MRAM[771][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8282_ (.D(_0378_),
    .CLK(net314),
    .Q(\mod.Data_Mem.F_M.MRAM[771][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8283_ (.D(_0379_),
    .CLK(net296),
    .Q(\mod.Data_Mem.F_M.MRAM[771][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8284_ (.D(_0380_),
    .CLK(net110),
    .Q(\mod.Data_Mem.F_M.MRAM[771][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8285_ (.D(_0381_),
    .CLK(net124),
    .Q(\mod.Data_Mem.F_M.MRAM[771][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8286_ (.D(_0382_),
    .CLK(net121),
    .Q(\mod.Data_Mem.F_M.MRAM[771][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8287_ (.D(_0383_),
    .CLK(net121),
    .Q(\mod.Data_Mem.F_M.MRAM[771][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8288_ (.D(_0384_),
    .CLK(net150),
    .Q(\mod.Data_Mem.F_M.MRAM[772][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8289_ (.D(_0385_),
    .CLK(net184),
    .Q(\mod.Data_Mem.F_M.MRAM[772][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8290_ (.D(_0386_),
    .CLK(net185),
    .Q(\mod.Data_Mem.F_M.MRAM[772][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8291_ (.D(_0387_),
    .CLK(net139),
    .Q(\mod.Data_Mem.F_M.MRAM[772][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8292_ (.D(_0388_),
    .CLK(net95),
    .Q(\mod.Data_Mem.F_M.MRAM[772][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8293_ (.D(_0389_),
    .CLK(net143),
    .Q(\mod.Data_Mem.F_M.MRAM[772][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8294_ (.D(_0390_),
    .CLK(net91),
    .Q(\mod.Data_Mem.F_M.MRAM[772][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8295_ (.D(_0391_),
    .CLK(net83),
    .Q(\mod.Data_Mem.F_M.MRAM[772][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8296_ (.D(_0392_),
    .CLK(net151),
    .Q(\mod.Data_Mem.F_M.MRAM[773][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8297_ (.D(_0393_),
    .CLK(net185),
    .Q(\mod.Data_Mem.F_M.MRAM[773][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8298_ (.D(_0394_),
    .CLK(net196),
    .Q(\mod.Data_Mem.F_M.MRAM[773][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8299_ (.D(_0395_),
    .CLK(net143),
    .Q(\mod.Data_Mem.F_M.MRAM[773][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8300_ (.D(_0396_),
    .CLK(net95),
    .Q(\mod.Data_Mem.F_M.MRAM[773][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8301_ (.D(_0397_),
    .CLK(net142),
    .Q(\mod.Data_Mem.F_M.MRAM[773][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8302_ (.D(_0398_),
    .CLK(net86),
    .Q(\mod.Data_Mem.F_M.MRAM[773][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8303_ (.D(_0399_),
    .CLK(net83),
    .Q(\mod.Data_Mem.F_M.MRAM[773][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8304_ (.D(_0400_),
    .CLK(net160),
    .Q(\mod.Data_Mem.F_M.MRAM[774][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8305_ (.D(_0401_),
    .CLK(net170),
    .Q(\mod.Data_Mem.F_M.MRAM[774][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8306_ (.D(_0402_),
    .CLK(net190),
    .Q(\mod.Data_Mem.F_M.MRAM[774][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8307_ (.D(_0403_),
    .CLK(net161),
    .Q(\mod.Data_Mem.F_M.MRAM[774][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8308_ (.D(_0404_),
    .CLK(net79),
    .Q(\mod.Data_Mem.F_M.MRAM[774][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8309_ (.D(_0405_),
    .CLK(net158),
    .Q(\mod.Data_Mem.F_M.MRAM[774][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8310_ (.D(_0406_),
    .CLK(net85),
    .Q(\mod.Data_Mem.F_M.MRAM[774][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8311_ (.D(_0407_),
    .CLK(net79),
    .Q(\mod.Data_Mem.F_M.MRAM[774][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8312_ (.D(_0408_),
    .CLK(net158),
    .Q(\mod.Data_Mem.F_M.MRAM[775][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8313_ (.D(_0409_),
    .CLK(net190),
    .Q(\mod.Data_Mem.F_M.MRAM[775][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8314_ (.D(_0410_),
    .CLK(net191),
    .Q(\mod.Data_Mem.F_M.MRAM[775][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8315_ (.D(_0411_),
    .CLK(net142),
    .Q(\mod.Data_Mem.F_M.MRAM[775][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8316_ (.D(_0412_),
    .CLK(net83),
    .Q(\mod.Data_Mem.F_M.MRAM[775][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8317_ (.D(_0413_),
    .CLK(net158),
    .Q(\mod.Data_Mem.F_M.MRAM[775][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8318_ (.D(_0414_),
    .CLK(net85),
    .Q(\mod.Data_Mem.F_M.MRAM[775][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8319_ (.D(_0415_),
    .CLK(net79),
    .Q(\mod.Data_Mem.F_M.MRAM[775][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8320_ (.D(_0416_),
    .CLK(net375),
    .Q(\mod.Data_Mem.F_M.MRAM[776][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8321_ (.D(_0417_),
    .CLK(net303),
    .Q(\mod.Data_Mem.F_M.MRAM[776][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8322_ (.D(_0418_),
    .CLK(net370),
    .Q(\mod.Data_Mem.F_M.MRAM[776][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8323_ (.D(_0419_),
    .CLK(net370),
    .Q(\mod.Data_Mem.F_M.MRAM[776][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8324_ (.D(_0420_),
    .CLK(net205),
    .Q(\mod.Data_Mem.F_M.MRAM[776][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8325_ (.D(_0421_),
    .CLK(net166),
    .Q(\mod.Data_Mem.F_M.MRAM[776][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8326_ (.D(_0422_),
    .CLK(net382),
    .Q(\mod.Data_Mem.F_M.MRAM[776][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8327_ (.D(_0423_),
    .CLK(net192),
    .Q(\mod.Data_Mem.F_M.MRAM[776][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8328_ (.D(_0424_),
    .CLK(net197),
    .Q(\mod.Data_Mem.F_M.MRAM[777][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8329_ (.D(_0425_),
    .CLK(net371),
    .Q(\mod.Data_Mem.F_M.MRAM[777][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8330_ (.D(_0426_),
    .CLK(net169),
    .Q(\mod.Data_Mem.F_M.MRAM[777][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8331_ (.D(_0427_),
    .CLK(net172),
    .Q(\mod.Data_Mem.F_M.MRAM[777][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8332_ (.D(_0428_),
    .CLK(net210),
    .Q(\mod.Data_Mem.F_M.MRAM[777][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8333_ (.D(_0429_),
    .CLK(net308),
    .Q(\mod.Data_Mem.F_M.MRAM[777][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8334_ (.D(_0430_),
    .CLK(net313),
    .Q(\mod.Data_Mem.F_M.MRAM[777][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8335_ (.D(_0431_),
    .CLK(net370),
    .Q(\mod.Data_Mem.F_M.MRAM[777][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8336_ (.D(_0432_),
    .CLK(net155),
    .Q(\mod.Data_Mem.F_M.MRAM[778][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8337_ (.D(_0433_),
    .CLK(net211),
    .Q(\mod.Data_Mem.F_M.MRAM[778][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8338_ (.D(_0434_),
    .CLK(net375),
    .Q(\mod.Data_Mem.F_M.MRAM[778][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8339_ (.D(_0435_),
    .CLK(net308),
    .Q(\mod.Data_Mem.F_M.MRAM[778][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8340_ (.D(_0436_),
    .CLK(net205),
    .Q(\mod.Data_Mem.F_M.MRAM[778][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8341_ (.D(_0437_),
    .CLK(net371),
    .Q(\mod.Data_Mem.F_M.MRAM[778][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8342_ (.D(_0438_),
    .CLK(net385),
    .Q(\mod.Data_Mem.F_M.MRAM[778][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8343_ (.D(_0439_),
    .CLK(net156),
    .Q(\mod.Data_Mem.F_M.MRAM[778][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8344_ (.D(_0440_),
    .CLK(net312),
    .Q(\mod.Data_Mem.F_M.MRAM[780][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8345_ (.D(_0441_),
    .CLK(net315),
    .Q(\mod.Data_Mem.F_M.MRAM[780][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8346_ (.D(_0442_),
    .CLK(net314),
    .Q(\mod.Data_Mem.F_M.MRAM[780][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8347_ (.D(_0443_),
    .CLK(net254),
    .Q(\mod.Data_Mem.F_M.MRAM[780][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8348_ (.D(_0444_),
    .CLK(net230),
    .Q(\mod.Data_Mem.F_M.MRAM[780][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8349_ (.D(_0445_),
    .CLK(net230),
    .Q(\mod.Data_Mem.F_M.MRAM[780][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8350_ (.D(_0446_),
    .CLK(net229),
    .Q(\mod.Data_Mem.F_M.MRAM[780][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8351_ (.D(_0447_),
    .CLK(net229),
    .Q(\mod.Data_Mem.F_M.MRAM[780][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8352_ (.D(_0448_),
    .CLK(net291),
    .Q(\mod.Data_Mem.F_M.MRAM[781][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8353_ (.D(_0449_),
    .CLK(net293),
    .Q(\mod.Data_Mem.F_M.MRAM[781][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8354_ (.D(_0450_),
    .CLK(net292),
    .Q(\mod.Data_Mem.F_M.MRAM[781][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8355_ (.D(_0451_),
    .CLK(net254),
    .Q(\mod.Data_Mem.F_M.MRAM[781][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8356_ (.D(_0452_),
    .CLK(net221),
    .Q(\mod.Data_Mem.F_M.MRAM[781][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8357_ (.D(_0453_),
    .CLK(net230),
    .Q(\mod.Data_Mem.F_M.MRAM[781][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8358_ (.D(_0454_),
    .CLK(net222),
    .Q(\mod.Data_Mem.F_M.MRAM[781][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8359_ (.D(_0455_),
    .CLK(net226),
    .Q(\mod.Data_Mem.F_M.MRAM[781][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8360_ (.D(_0456_),
    .CLK(net287),
    .Q(\mod.Data_Mem.F_M.MRAM[782][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8361_ (.D(_0457_),
    .CLK(net293),
    .Q(\mod.Data_Mem.F_M.MRAM[782][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8362_ (.D(_0458_),
    .CLK(net292),
    .Q(\mod.Data_Mem.F_M.MRAM[782][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8363_ (.D(_0459_),
    .CLK(net254),
    .Q(\mod.Data_Mem.F_M.MRAM[782][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8364_ (.D(_0460_),
    .CLK(net221),
    .Q(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8365_ (.D(_0461_),
    .CLK(net229),
    .Q(\mod.Data_Mem.F_M.MRAM[782][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8366_ (.D(_0462_),
    .CLK(net221),
    .Q(\mod.Data_Mem.F_M.MRAM[782][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8367_ (.D(_0463_),
    .CLK(net221),
    .Q(\mod.Data_Mem.F_M.MRAM[782][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8368_ (.D(_0464_),
    .CLK(net287),
    .Q(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8369_ (.D(_0465_),
    .CLK(net291),
    .Q(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8370_ (.D(_0466_),
    .CLK(net292),
    .Q(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8371_ (.D(_0467_),
    .CLK(net255),
    .Q(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8372_ (.D(_0468_),
    .CLK(net229),
    .Q(\mod.Data_Mem.F_M.MRAM[783][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8373_ (.D(_0469_),
    .CLK(net127),
    .Q(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8374_ (.D(_0470_),
    .CLK(net119),
    .Q(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8375_ (.D(_0471_),
    .CLK(net119),
    .Q(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8376_ (.D(_0472_),
    .CLK(net215),
    .Q(\mod.Data_Mem.F_M.MRAM[784][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8377_ (.D(_0473_),
    .CLK(net316),
    .Q(\mod.Data_Mem.F_M.MRAM[784][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8378_ (.D(_0474_),
    .CLK(net316),
    .Q(\mod.Data_Mem.F_M.MRAM[784][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8379_ (.D(_0475_),
    .CLK(net180),
    .Q(\mod.Data_Mem.F_M.MRAM[784][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8380_ (.D(_0476_),
    .CLK(net120),
    .Q(\mod.Data_Mem.F_M.MRAM[784][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8381_ (.D(_0477_),
    .CLK(net110),
    .Q(\mod.Data_Mem.F_M.MRAM[784][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8382_ (.D(_0478_),
    .CLK(net116),
    .Q(\mod.Data_Mem.F_M.MRAM[784][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8383_ (.D(_0479_),
    .CLK(net117),
    .Q(\mod.Data_Mem.F_M.MRAM[784][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8384_ (.D(_0480_),
    .CLK(net180),
    .Q(\mod.Data_Mem.F_M.MRAM[785][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8385_ (.D(_0481_),
    .CLK(net181),
    .Q(\mod.Data_Mem.F_M.MRAM[785][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8386_ (.D(_0482_),
    .CLK(net181),
    .Q(\mod.Data_Mem.F_M.MRAM[785][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8387_ (.D(_0483_),
    .CLK(net180),
    .Q(\mod.Data_Mem.F_M.MRAM[785][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8388_ (.D(_0484_),
    .CLK(net104),
    .Q(\mod.Data_Mem.F_M.MRAM[785][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8389_ (.D(_0485_),
    .CLK(net105),
    .Q(\mod.Data_Mem.F_M.MRAM[785][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8390_ (.D(_0486_),
    .CLK(net74),
    .Q(\mod.Data_Mem.F_M.MRAM[785][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8391_ (.D(_0487_),
    .CLK(net77),
    .Q(\mod.Data_Mem.F_M.MRAM[785][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8392_ (.D(_0488_),
    .CLK(net179),
    .Q(\mod.Data_Mem.F_M.MRAM[786][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8393_ (.D(_0489_),
    .CLK(net201),
    .Q(\mod.Data_Mem.F_M.MRAM[786][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8394_ (.D(_0490_),
    .CLK(net201),
    .Q(\mod.Data_Mem.F_M.MRAM[786][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8395_ (.D(_0491_),
    .CLK(net179),
    .Q(\mod.Data_Mem.F_M.MRAM[786][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8396_ (.D(_0492_),
    .CLK(net104),
    .Q(\mod.Data_Mem.F_M.MRAM[786][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8397_ (.D(_0493_),
    .CLK(net105),
    .Q(\mod.Data_Mem.F_M.MRAM[786][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8398_ (.D(_0494_),
    .CLK(net104),
    .Q(\mod.Data_Mem.F_M.MRAM[786][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8399_ (.D(_0495_),
    .CLK(net104),
    .Q(\mod.Data_Mem.F_M.MRAM[786][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8400_ (.D(_0496_),
    .CLK(net179),
    .Q(\mod.Data_Mem.F_M.MRAM[787][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8401_ (.D(_0497_),
    .CLK(net182),
    .Q(\mod.Data_Mem.F_M.MRAM[787][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8402_ (.D(_0498_),
    .CLK(net182),
    .Q(\mod.Data_Mem.F_M.MRAM[787][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8403_ (.D(_0499_),
    .CLK(net179),
    .Q(\mod.Data_Mem.F_M.MRAM[787][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8404_ (.D(_0500_),
    .CLK(net97),
    .Q(\mod.Data_Mem.F_M.MRAM[787][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8405_ (.D(_0501_),
    .CLK(net105),
    .Q(\mod.Data_Mem.F_M.MRAM[787][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8406_ (.D(_0502_),
    .CLK(net97),
    .Q(\mod.Data_Mem.F_M.MRAM[787][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8407_ (.D(_0503_),
    .CLK(net97),
    .Q(\mod.Data_Mem.F_M.MRAM[787][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8408_ (.D(_0504_),
    .CLK(net140),
    .Q(\mod.Data_Mem.F_M.MRAM[788][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8409_ (.D(_0505_),
    .CLK(net160),
    .Q(\mod.Data_Mem.F_M.MRAM[788][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8410_ (.D(_0506_),
    .CLK(net190),
    .Q(\mod.Data_Mem.F_M.MRAM[788][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8411_ (.D(_0507_),
    .CLK(net142),
    .Q(\mod.Data_Mem.F_M.MRAM[788][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8412_ (.D(_0508_),
    .CLK(net85),
    .Q(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8413_ (.D(_0509_),
    .CLK(net139),
    .Q(\mod.Data_Mem.F_M.MRAM[788][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8414_ (.D(_0510_),
    .CLK(net87),
    .Q(\mod.Data_Mem.F_M.MRAM[788][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8415_ (.D(_0511_),
    .CLK(net88),
    .Q(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8416_ (.D(_0512_),
    .CLK(net149),
    .Q(\mod.Data_Mem.F_M.MRAM[790][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8417_ (.D(_0513_),
    .CLK(net150),
    .Q(\mod.Data_Mem.F_M.MRAM[790][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8418_ (.D(_0514_),
    .CLK(net188),
    .Q(\mod.Data_Mem.F_M.MRAM[790][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8419_ (.D(_0515_),
    .CLK(net138),
    .Q(\mod.Data_Mem.F_M.MRAM[790][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8420_ (.D(_0516_),
    .CLK(net86),
    .Q(\mod.Data_Mem.F_M.MRAM[790][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8421_ (.D(_0517_),
    .CLK(net162),
    .Q(\mod.Data_Mem.F_M.MRAM[790][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8422_ (.D(_0518_),
    .CLK(net86),
    .Q(\mod.Data_Mem.F_M.MRAM[790][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8423_ (.D(_0519_),
    .CLK(net92),
    .Q(\mod.Data_Mem.F_M.MRAM[790][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8424_ (.D(_0520_),
    .CLK(net147),
    .Q(\mod.Data_Mem.F_M.MRAM[791][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8425_ (.D(_0521_),
    .CLK(net150),
    .Q(\mod.Data_Mem.F_M.MRAM[791][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8426_ (.D(_0522_),
    .CLK(net188),
    .Q(\mod.Data_Mem.F_M.MRAM[791][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8427_ (.D(_0523_),
    .CLK(net138),
    .Q(\mod.Data_Mem.F_M.MRAM[791][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8428_ (.D(_0524_),
    .CLK(net87),
    .Q(\mod.Data_Mem.F_M.MRAM[791][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8429_ (.D(_0525_),
    .CLK(net162),
    .Q(\mod.Data_Mem.F_M.MRAM[791][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8430_ (.D(_0526_),
    .CLK(net91),
    .Q(\mod.Data_Mem.F_M.MRAM[791][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8431_ (.D(_0527_),
    .CLK(net90),
    .Q(\mod.Data_Mem.F_M.MRAM[791][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8432_ (.D(_0528_),
    .CLK(net192),
    .Q(\mod.Data_Mem.F_M.MRAM[792][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8433_ (.D(_0529_),
    .CLK(net193),
    .Q(\mod.Data_Mem.F_M.MRAM[792][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8434_ (.D(_0530_),
    .CLK(net323),
    .Q(\mod.Data_Mem.F_M.MRAM[792][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8435_ (.D(_0531_),
    .CLK(net377),
    .Q(\mod.Data_Mem.F_M.MRAM[792][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8436_ (.D(_0532_),
    .CLK(net155),
    .Q(\mod.Data_Mem.F_M.MRAM[792][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8437_ (.D(_0533_),
    .CLK(net192),
    .Q(\mod.Data_Mem.F_M.MRAM[792][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8438_ (.D(_0534_),
    .CLK(net379),
    .Q(\mod.Data_Mem.F_M.MRAM[792][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8439_ (.D(_0535_),
    .CLK(net373),
    .Q(\mod.Data_Mem.F_M.MRAM[792][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8440_ (.D(_0536_),
    .CLK(net320),
    .Q(\mod.Data_Mem.F_M.MRAM[793][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8441_ (.D(_0537_),
    .CLK(net198),
    .Q(\mod.Data_Mem.F_M.MRAM[793][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8442_ (.D(_0538_),
    .CLK(net156),
    .Q(\mod.Data_Mem.F_M.MRAM[793][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8443_ (.D(_0539_),
    .CLK(net166),
    .Q(\mod.Data_Mem.F_M.MRAM[793][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8444_ (.D(_0540_),
    .CLK(net192),
    .Q(\mod.Data_Mem.F_M.MRAM[793][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8445_ (.D(_0541_),
    .CLK(net377),
    .Q(\mod.Data_Mem.F_M.MRAM[793][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8446_ (.D(_0542_),
    .CLK(net373),
    .Q(\mod.Data_Mem.F_M.MRAM[793][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8447_ (.D(_0543_),
    .CLK(net342),
    .Q(\mod.Data_Mem.F_M.MRAM[793][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8448_ (.D(_0544_),
    .CLK(net372),
    .Q(\mod.Data_Mem.F_M.MRAM[794][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8449_ (.D(_0545_),
    .CLK(net376),
    .Q(\mod.Data_Mem.F_M.MRAM[794][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8450_ (.D(_0546_),
    .CLK(net167),
    .Q(\mod.Data_Mem.F_M.MRAM[794][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8451_ (.D(_0547_),
    .CLK(net377),
    .Q(\mod.Data_Mem.F_M.MRAM[794][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8452_ (.D(_0548_),
    .CLK(net375),
    .Q(\mod.Data_Mem.F_M.MRAM[794][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8453_ (.D(_0549_),
    .CLK(net315),
    .Q(\mod.Data_Mem.F_M.MRAM[794][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8454_ (.D(_0550_),
    .CLK(net168),
    .Q(\mod.Data_Mem.F_M.MRAM[794][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8455_ (.D(_0551_),
    .CLK(net369),
    .Q(\mod.Data_Mem.F_M.MRAM[794][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8456_ (.D(_0552_),
    .CLK(net317),
    .Q(\mod.Data_Mem.F_M.MRAM[795][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8457_ (.D(_0553_),
    .CLK(net368),
    .Q(\mod.Data_Mem.F_M.MRAM[795][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8458_ (.D(_0554_),
    .CLK(net323),
    .Q(\mod.Data_Mem.F_M.MRAM[795][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8459_ (.D(_0555_),
    .CLK(net387),
    .Q(\mod.Data_Mem.F_M.MRAM[795][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8460_ (.D(_0556_),
    .CLK(net173),
    .Q(\mod.Data_Mem.F_M.MRAM[795][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8461_ (.D(_0557_),
    .CLK(net157),
    .Q(\mod.Data_Mem.F_M.MRAM[795][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8462_ (.D(_0558_),
    .CLK(net384),
    .Q(\mod.Data_Mem.F_M.MRAM[795][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8463_ (.D(_0559_),
    .CLK(net321),
    .Q(\mod.Data_Mem.F_M.MRAM[795][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8464_ (.D(_0560_),
    .CLK(net287),
    .Q(\mod.Data_Mem.F_M.MRAM[796][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8465_ (.D(_0561_),
    .CLK(net291),
    .Q(\mod.Data_Mem.F_M.MRAM[796][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8466_ (.D(_0562_),
    .CLK(net292),
    .Q(\mod.Data_Mem.F_M.MRAM[796][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8467_ (.D(_0563_),
    .CLK(net288),
    .Q(\mod.Data_Mem.F_M.MRAM[796][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8468_ (.D(_0564_),
    .CLK(net236),
    .Q(\mod.Data_Mem.F_M.MRAM[796][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8469_ (.D(_0565_),
    .CLK(net235),
    .Q(\mod.Data_Mem.F_M.MRAM[796][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8470_ (.D(_0566_),
    .CLK(net237),
    .Q(\mod.Data_Mem.F_M.MRAM[796][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8471_ (.D(_0567_),
    .CLK(net238),
    .Q(\mod.Data_Mem.F_M.MRAM[796][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8472_ (.D(_0568_),
    .CLK(net287),
    .Q(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8473_ (.D(_0569_),
    .CLK(net291),
    .Q(\mod.Data_Mem.F_M.MRAM[797][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8474_ (.D(_0570_),
    .CLK(net293),
    .Q(\mod.Data_Mem.F_M.MRAM[797][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8475_ (.D(_0571_),
    .CLK(net288),
    .Q(\mod.Data_Mem.F_M.MRAM[797][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8476_ (.D(_0572_),
    .CLK(net236),
    .Q(\mod.Data_Mem.F_M.MRAM[797][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8477_ (.D(_0573_),
    .CLK(net235),
    .Q(\mod.Data_Mem.F_M.MRAM[797][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8478_ (.D(_0574_),
    .CLK(net237),
    .Q(\mod.Data_Mem.F_M.MRAM[797][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8479_ (.D(_0575_),
    .CLK(net238),
    .Q(\mod.Data_Mem.F_M.MRAM[797][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8480_ (.D(_0576_),
    .CLK(net289),
    .Q(\mod.Data_Mem.F_M.MRAM[798][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8481_ (.D(_0577_),
    .CLK(net294),
    .Q(\mod.Data_Mem.F_M.MRAM[798][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8482_ (.D(_0578_),
    .CLK(net341),
    .Q(\mod.Data_Mem.F_M.MRAM[798][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8483_ (.D(_0579_),
    .CLK(net256),
    .Q(\mod.Data_Mem.F_M.MRAM[798][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8484_ (.D(_0580_),
    .CLK(net101),
    .Q(\mod.Data_Mem.F_M.MRAM[798][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8485_ (.D(_0581_),
    .CLK(net110),
    .Q(\mod.Data_Mem.F_M.MRAM[798][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8486_ (.D(_0582_),
    .CLK(net102),
    .Q(\mod.Data_Mem.F_M.MRAM[798][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8487_ (.D(_0583_),
    .CLK(net102),
    .Q(\mod.Data_Mem.F_M.MRAM[798][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8488_ (.D(_0584_),
    .CLK(net164),
    .Q(\mod.Data_Mem.F_M.MRAM[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8489_ (.D(_0585_),
    .CLK(net140),
    .Q(\mod.Data_Mem.F_M.MRAM[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8490_ (.D(_0586_),
    .CLK(net145),
    .Q(\mod.Data_Mem.F_M.MRAM[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8491_ (.D(_0587_),
    .CLK(net386),
    .Q(\mod.Data_Mem.F_M.MRAM[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8492_ (.D(_0588_),
    .CLK(net84),
    .Q(\mod.Data_Mem.F_M.MRAM[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8493_ (.D(_0589_),
    .CLK(net160),
    .Q(\mod.Data_Mem.F_M.MRAM[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8494_ (.D(_0590_),
    .CLK(net80),
    .Q(\mod.Data_Mem.F_M.MRAM[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8495_ (.D(_0591_),
    .CLK(net72),
    .Q(\mod.Data_Mem.F_M.MRAM[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8496_ (.D(_0000_),
    .CLK(net268),
    .Q(\mod.Data_Mem.F_M.out_data[72] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8497_ (.D(_0001_),
    .CLK(net268),
    .Q(\mod.Data_Mem.F_M.out_data[73] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8498_ (.D(_0002_),
    .CLK(net339),
    .Q(\mod.Data_Mem.F_M.out_data[74] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8499_ (.D(_0003_),
    .CLK(net265),
    .Q(\mod.Data_Mem.F_M.out_data[75] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8500_ (.D(_0004_),
    .CLK(net246),
    .Q(\mod.Data_Mem.F_M.out_data[76] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8501_ (.D(_0005_),
    .CLK(net265),
    .Q(\mod.Data_Mem.F_M.out_data[77] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8502_ (.D(_0006_),
    .CLK(net264),
    .Q(\mod.Data_Mem.F_M.out_data[78] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8503_ (.D(_0007_),
    .CLK(net246),
    .Q(\mod.Data_Mem.F_M.out_data[79] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8504_ (.D(_0008_),
    .CLK(net349),
    .Q(\mod.Data_Mem.F_M.out_data[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8505_ (.D(_0009_),
    .CLK(net335),
    .Q(\mod.Data_Mem.F_M.out_data[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8506_ (.D(_0010_),
    .CLK(net348),
    .Q(\mod.Data_Mem.F_M.out_data[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8507_ (.D(_0011_),
    .CLK(net345),
    .Q(\mod.Data_Mem.F_M.out_data[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8508_ (.D(net573),
    .CLK(net359),
    .Q(\mod.Data_Mem.F_M.out_data[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8509_ (.D(net572),
    .CLK(net357),
    .Q(\mod.Data_Mem.F_M.out_data[69] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8510_ (.D(net571),
    .CLK(net383),
    .Q(\mod.Data_Mem.F_M.out_data[70] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8511_ (.D(net570),
    .CLK(net358),
    .Q(\mod.Data_Mem.F_M.out_data[71] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8512_ (.D(_0016_),
    .CLK(net340),
    .Q(\mod.Data_Mem.F_M.out_data[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8513_ (.D(_0017_),
    .CLK(net330),
    .Q(\mod.Data_Mem.F_M.out_data[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8514_ (.D(_0018_),
    .CLK(net331),
    .Q(\mod.Data_Mem.F_M.out_data[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8515_ (.D(_0019_),
    .CLK(net355),
    .Q(\mod.Data_Mem.F_M.out_data[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8516_ (.D(net569),
    .CLK(net359),
    .Q(\mod.Data_Mem.F_M.out_data[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8517_ (.D(net568),
    .CLK(net362),
    .Q(\mod.Data_Mem.F_M.out_data[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8518_ (.D(net567),
    .CLK(net362),
    .Q(\mod.Data_Mem.F_M.out_data[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8519_ (.D(net566),
    .CLK(net361),
    .Q(\mod.Data_Mem.F_M.out_data[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8520_ (.D(_0024_),
    .CLK(net350),
    .Q(\mod.Data_Mem.F_M.out_data[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8521_ (.D(_0025_),
    .CLK(net332),
    .Q(\mod.Data_Mem.F_M.out_data[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8522_ (.D(_0026_),
    .CLK(net340),
    .Q(\mod.Data_Mem.F_M.out_data[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8523_ (.D(_0027_),
    .CLK(net355),
    .Q(\mod.Data_Mem.F_M.out_data[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8524_ (.D(net565),
    .CLK(net357),
    .Q(\mod.Data_Mem.F_M.out_data[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8525_ (.D(net564),
    .CLK(net357),
    .Q(\mod.Data_Mem.F_M.out_data[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8526_ (.D(net563),
    .CLK(net363),
    .Q(\mod.Data_Mem.F_M.out_data[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8527_ (.D(net562),
    .CLK(net363),
    .Q(\mod.Data_Mem.F_M.out_data[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8528_ (.D(_0032_),
    .CLK(net330),
    .Q(\mod.Data_Mem.F_M.out_data[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8529_ (.D(_0033_),
    .CLK(net332),
    .Q(\mod.Data_Mem.F_M.out_data[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8530_ (.D(_0034_),
    .CLK(net288),
    .Q(\mod.Data_Mem.F_M.out_data[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8531_ (.D(_0035_),
    .CLK(net328),
    .Q(\mod.Data_Mem.F_M.out_data[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8532_ (.D(_0036_),
    .CLK(net252),
    .Q(\mod.Data_Mem.F_M.out_data[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8533_ (.D(_0037_),
    .CLK(net277),
    .Q(\mod.Data_Mem.F_M.out_data[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8534_ (.D(_0038_),
    .CLK(net253),
    .Q(\mod.Data_Mem.F_M.out_data[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8535_ (.D(_0039_),
    .CLK(net254),
    .Q(\mod.Data_Mem.F_M.out_data[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8536_ (.D(_0040_),
    .CLK(net330),
    .Q(\mod.Data_Mem.F_M.out_data[32] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8537_ (.D(_0041_),
    .CLK(net344),
    .Q(\mod.Data_Mem.F_M.out_data[33] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8538_ (.D(_0042_),
    .CLK(net346),
    .Q(\mod.Data_Mem.F_M.out_data[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8539_ (.D(_0043_),
    .CLK(net277),
    .Q(\mod.Data_Mem.F_M.out_data[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8540_ (.D(_0044_),
    .CLK(net269),
    .Q(\mod.Data_Mem.F_M.out_data[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8541_ (.D(_0045_),
    .CLK(net271),
    .Q(\mod.Data_Mem.F_M.out_data[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8542_ (.D(_0046_),
    .CLK(net253),
    .Q(\mod.Data_Mem.F_M.out_data[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8543_ (.D(_0047_),
    .CLK(net251),
    .Q(\mod.Data_Mem.F_M.out_data[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8544_ (.D(_0048_),
    .CLK(net327),
    .Q(\mod.Data_Mem.F_M.out_data[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8545_ (.D(_0049_),
    .CLK(net327),
    .Q(\mod.Data_Mem.F_M.out_data[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8546_ (.D(_0050_),
    .CLK(net331),
    .Q(\mod.Data_Mem.F_M.out_data[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8547_ (.D(_0051_),
    .CLK(net327),
    .Q(\mod.Data_Mem.F_M.out_data[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8548_ (.D(_0052_),
    .CLK(net252),
    .Q(\mod.Data_Mem.F_M.out_data[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8549_ (.D(_0053_),
    .CLK(net277),
    .Q(\mod.Data_Mem.F_M.out_data[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8550_ (.D(_0054_),
    .CLK(net252),
    .Q(\mod.Data_Mem.F_M.out_data[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8551_ (.D(_0055_),
    .CLK(net251),
    .Q(\mod.Data_Mem.F_M.out_data[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8552_ (.D(_0056_),
    .CLK(net256),
    .Q(\mod.Data_Mem.F_M.out_data[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8553_ (.D(_0057_),
    .CLK(net342),
    .Q(\mod.Data_Mem.F_M.out_data[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8554_ (.D(_0058_),
    .CLK(net342),
    .Q(\mod.Data_Mem.F_M.out_data[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8555_ (.D(_0059_),
    .CLK(net328),
    .Q(\mod.Data_Mem.F_M.out_data[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8556_ (.D(_0060_),
    .CLK(net277),
    .Q(\mod.Data_Mem.F_M.out_data[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8557_ (.D(_0061_),
    .CLK(net280),
    .Q(\mod.Data_Mem.F_M.out_data[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8558_ (.D(_0062_),
    .CLK(net275),
    .Q(\mod.Data_Mem.F_M.out_data[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8559_ (.D(_0063_),
    .CLK(net275),
    .Q(\mod.Data_Mem.F_M.out_data[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8560_ (.D(_0064_),
    .CLK(net339),
    .Q(\mod.Data_Mem.F_M.out_data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8561_ (.D(_0065_),
    .CLK(net340),
    .Q(\mod.Data_Mem.F_M.out_data[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8562_ (.D(_0066_),
    .CLK(net347),
    .Q(\mod.Data_Mem.F_M.out_data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8563_ (.D(_0067_),
    .CLK(net337),
    .Q(\mod.Data_Mem.F_M.out_data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8564_ (.D(_0068_),
    .CLK(net248),
    .Q(\mod.Data_Mem.F_M.out_data[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8565_ (.D(_0069_),
    .CLK(net247),
    .Q(\mod.Data_Mem.F_M.out_data[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8566_ (.D(_0070_),
    .CLK(net248),
    .Q(\mod.Data_Mem.F_M.out_data[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8567_ (.D(_0071_),
    .CLK(net247),
    .Q(\mod.Data_Mem.F_M.out_data[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8568_ (.D(_0072_),
    .CLK(net340),
    .Q(\mod.Data_Mem.F_M.out_data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8569_ (.D(_0073_),
    .CLK(net349),
    .Q(\mod.Data_Mem.F_M.out_data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8570_ (.D(_0074_),
    .CLK(net349),
    .Q(\mod.Data_Mem.F_M.out_data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8571_ (.D(_0075_),
    .CLK(net334),
    .Q(\mod.Data_Mem.F_M.out_data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8572_ (.D(_0076_),
    .CLK(net247),
    .Q(\mod.Data_Mem.F_M.out_data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8573_ (.D(_0077_),
    .CLK(net282),
    .Q(\mod.Data_Mem.F_M.out_data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8574_ (.D(_0078_),
    .CLK(net264),
    .Q(\mod.Data_Mem.F_M.out_data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8575_ (.D(_0079_),
    .CLK(net245),
    .Q(\mod.Data_Mem.F_M.out_data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8576_ (.D(_0592_),
    .CLK(net263),
    .Q(\mod.Instr_Mem.instruction[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8577_ (.D(_0593_),
    .CLK(net117),
    .Q(\mod.Instr_Mem.instruction[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8578_ (.D(_0594_),
    .CLK(net263),
    .Q(\mod.Instr_Mem.instruction[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8579_ (.D(_0595_),
    .CLK(net218),
    .Q(\mod.Instr_Mem.instruction[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8580_ (.D(_0596_),
    .CLK(net119),
    .Q(\mod.Instr_Mem.instruction[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8581_ (.D(_0597_),
    .CLK(net218),
    .Q(\mod.Instr_Mem.instruction[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8582_ (.D(_0598_),
    .CLK(net100),
    .Q(\mod.Instr_Mem.instruction[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8583_ (.D(_0599_),
    .CLK(net101),
    .Q(\mod.Instr_Mem.instruction[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8584_ (.D(_0600_),
    .CLK(net171),
    .Q(\mod.Data_Mem.F_M.MRAM[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8585_ (.D(_0601_),
    .CLK(net168),
    .Q(\mod.Data_Mem.F_M.MRAM[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8586_ (.D(_0602_),
    .CLK(net378),
    .Q(\mod.Data_Mem.F_M.MRAM[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8587_ (.D(_0603_),
    .CLK(net371),
    .Q(\mod.Data_Mem.F_M.MRAM[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8588_ (.D(_0604_),
    .CLK(net197),
    .Q(\mod.Data_Mem.F_M.MRAM[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8589_ (.D(_0605_),
    .CLK(net167),
    .Q(\mod.Data_Mem.F_M.MRAM[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8590_ (.D(_0606_),
    .CLK(net193),
    .Q(\mod.Data_Mem.F_M.MRAM[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8591_ (.D(_0607_),
    .CLK(net385),
    .Q(\mod.Data_Mem.F_M.MRAM[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8592_ (.D(_0608_),
    .CLK(net220),
    .Q(\mod.Instr_Mem.instruction[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8593_ (.D(_0609_),
    .CLK(net226),
    .Q(\mod.Instr_Mem.instruction[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8594_ (.D(_0610_),
    .CLK(net115),
    .Q(\mod.Instr_Mem.instruction[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8595_ (.D(_0611_),
    .CLK(net220),
    .Q(\mod.Instr_Mem.instruction[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__D (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_395 (.ZN(net395));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_396 (.ZN(net396));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_397 (.ZN(net397));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_398 (.ZN(net398));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_399 (.ZN(net399));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_400 (.ZN(net400));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_401 (.ZN(net401));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_402 (.ZN(net402));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_403 (.ZN(net403));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_404 (.ZN(net404));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_405 (.ZN(net405));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_406 (.ZN(net406));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_407 (.ZN(net407));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_408 (.ZN(net408));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_409 (.ZN(net409));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_410 (.ZN(net410));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_411 (.ZN(net411));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_412 (.ZN(net412));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_413 (.ZN(net413));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_414 (.ZN(net414));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_415 (.ZN(net415));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_416 (.ZN(net416));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_417 (.ZN(net417));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_418 (.ZN(net418));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_419 (.ZN(net419));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_420 (.ZN(net420));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_421 (.ZN(net421));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_422 (.ZN(net422));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_423 (.ZN(net423));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_424 (.ZN(net424));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_425 (.ZN(net425));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_426 (.ZN(net426));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_427 (.ZN(net427));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_428 (.ZN(net428));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_429 (.ZN(net429));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_430 (.ZN(net430));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_431 (.ZN(net431));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_432 (.ZN(net432));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_433 (.ZN(net433));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_434 (.ZN(net434));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_435 (.ZN(net435));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_436 (.ZN(net436));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_437 (.ZN(net437));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_438 (.ZN(net438));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_439 (.ZN(net439));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_440 (.ZN(net440));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_441 (.ZN(net441));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_442 (.ZN(net442));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_443 (.ZN(net443));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_444 (.ZN(net444));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_445 (.ZN(net445));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_446 (.ZN(net446));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_447 (.ZN(net447));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_448 (.ZN(net448));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_449 (.ZN(net449));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_450 (.ZN(net450));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_451 (.ZN(net451));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_452 (.ZN(net452));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_453 (.ZN(net453));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_454 (.ZN(net454));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_455 (.ZN(net455));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_456 (.ZN(net456));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_457 (.ZN(net457));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_458 (.ZN(net458));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_459 (.ZN(net459));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_460 (.ZN(net460));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_461 (.ZN(net461));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_462 (.ZN(net462));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_463 (.ZN(net463));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_464 (.ZN(net464));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_465 (.ZN(net465));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_466 (.ZN(net466));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_467 (.ZN(net467));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_468 (.ZN(net468));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_469 (.ZN(net469));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_470 (.ZN(net470));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_471 (.ZN(net471));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_472 (.ZN(net472));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_473 (.ZN(net473));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_474 (.ZN(net474));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_475 (.ZN(net475));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_476 (.ZN(net476));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_477 (.ZN(net477));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_478 (.ZN(net478));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_479 (.ZN(net479));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_480 (.ZN(net480));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_481 (.ZN(net481));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_482 (.ZN(net482));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_483 (.ZN(net483));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_484 (.ZN(net484));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_485 (.ZN(net485));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_486 (.ZN(net486));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_487 (.ZN(net487));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_488 (.ZN(net488));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_489 (.ZN(net489));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_490 (.ZN(net490));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_491 (.ZN(net491));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_492 (.ZN(net492));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_493 (.ZN(net493));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_494 (.ZN(net494));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_495 (.ZN(net495));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_496 (.ZN(net496));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_497 (.ZN(net497));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_498 (.ZN(net498));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_499 (.ZN(net499));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_500 (.ZN(net500));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_501 (.ZN(net501));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_502 (.ZN(net502));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_503 (.ZN(net503));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_504 (.ZN(net504));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_505 (.ZN(net505));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_506 (.ZN(net506));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_507 (.ZN(net507));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_508 (.ZN(net508));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_509 (.ZN(net509));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_510 (.ZN(net510));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_511 (.ZN(net511));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_512 (.ZN(net512));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_513 (.ZN(net513));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_514 (.ZN(net514));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_515 (.ZN(net515));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_516 (.ZN(net516));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_517 (.ZN(net517));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_518 (.ZN(net518));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_519 (.ZN(net519));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_520 (.ZN(net520));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_521 (.ZN(net521));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_522 (.ZN(net522));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_523 (.ZN(net523));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_524 (.ZN(net524));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_525 (.ZN(net525));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_526 (.ZN(net526));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_527 (.ZN(net527));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_528 (.ZN(net528));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_529 (.ZN(net529));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_530 (.ZN(net530));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_531 (.ZN(net531));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_532 (.ZN(net532));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_533 (.ZN(net533));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_534 (.ZN(net534));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_535 (.ZN(net535));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_536 (.ZN(net536));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_537 (.ZN(net537));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_538 (.ZN(net538));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_539 (.ZN(net539));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_540 (.ZN(net540));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_541 (.ZN(net541));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_542 (.ZN(net542));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_543 (.ZN(net543));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_544 (.ZN(net544));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_545 (.ZN(net545));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_546 (.ZN(net546));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_547 (.ZN(net547));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_548 (.ZN(net548));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_549 (.ZN(net549));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_550 (.ZN(net550));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_551 (.ZN(net551));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_552 (.ZN(net552));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_553 (.ZN(net553));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_554 (.ZN(net554));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_555 (.ZN(net555));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_556 (.ZN(net556));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_557 (.ZN(net557));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_558 (.ZN(net558));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_559 (.ZN(net559));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_560 (.ZN(net560));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_561 (.ZN(net561));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8527__562 (.ZN(net562));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8526__563 (.ZN(net563));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8525__564 (.ZN(net564));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8524__565 (.ZN(net565));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8519__566 (.ZN(net566));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8518__567 (.ZN(net567));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8517__568 (.ZN(net568));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8516__569 (.ZN(net569));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8511__570 (.ZN(net570));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8510__571 (.ZN(net571));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8509__572 (.ZN(net572));
 gf180mcu_fd_sc_mcu7t5v0__tiel _8508__573 (.ZN(net573));
 gf180mcu_fd_sc_mcu7t5v0__tieh _8194__574 (.Z(net574));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_in[8]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_in[9]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output3 (.I(net3),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output4 (.I(net4),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output5 (.I(net5),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output6 (.I(net6),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output8 (.I(net8),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output9 (.I(net9),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output10 (.I(net10),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout11 (.I(net13),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout12 (.I(net13),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout13 (.I(net15),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout14 (.I(net15),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout15 (.I(net24),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout16 (.I(net18),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout17 (.I(net18),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout18 (.I(net22),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout19 (.I(net22),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout20 (.I(net22),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout21 (.I(net22),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout22 (.I(net23),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout23 (.I(net24),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout24 (.I(net39),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout25 (.I(net38),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout26 (.I(net33),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout27 (.I(net33),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout28 (.I(net29),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout29 (.I(net31),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout30 (.I(net31),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout31 (.I(net32),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout32 (.I(net33),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout33 (.I(net37),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout34 (.I(net36),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout35 (.I(net36),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout36 (.I(net37),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout37 (.I(net38),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout38 (.I(net39),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout39 (.I(net69),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout40 (.I(net42),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout41 (.I(net42),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout42 (.I(net45),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout43 (.I(net45),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout44 (.I(net50),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout45 (.I(net50),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout47 (.I(net49),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net51),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout51 (.I(net68),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net53),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout53 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout54 (.I(net67),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout55 (.I(net56),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout56 (.I(net57),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout57 (.I(net66),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout58 (.I(net59),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout59 (.I(net65),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout60 (.I(net65),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout61 (.I(net62),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout62 (.I(net64),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout63 (.I(net65),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout64 (.I(net65),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout65 (.I(net66),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout68 (.I(net69),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout69 (.I(net2),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout70 (.I(net76),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout71 (.I(net72),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout72 (.I(net76),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout73 (.I(net75),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout74 (.I(net75),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout75 (.I(net76),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout76 (.I(net77),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout77 (.I(net96),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout78 (.I(net96),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout79 (.I(net80),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout80 (.I(net84),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout81 (.I(net82),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout82 (.I(net83),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout83 (.I(net84),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout84 (.I(net94),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout85 (.I(net87),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout86 (.I(net87),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout87 (.I(net90),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout89 (.I(net90),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout90 (.I(net93),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout91 (.I(net93),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout92 (.I(net93),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout93 (.I(net94),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout94 (.I(net95),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout95 (.I(net96),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout96 (.I(net137),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout97 (.I(net99),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout98 (.I(net99),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout99 (.I(net103),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout100 (.I(net101),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout101 (.I(net103),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout102 (.I(net103),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout103 (.I(net113),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout104 (.I(net108),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout105 (.I(net108),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout106 (.I(net108),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout107 (.I(net108),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout108 (.I(net112),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout109 (.I(net111),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout110 (.I(net112),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout111 (.I(net112),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout112 (.I(net113),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout113 (.I(net131),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout114 (.I(net115),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout115 (.I(net117),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout116 (.I(net117),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout117 (.I(net120),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout118 (.I(net119),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout119 (.I(net120),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout120 (.I(net130),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout121 (.I(net124),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout122 (.I(net123),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout123 (.I(net124),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout124 (.I(net129),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout125 (.I(net128),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout126 (.I(net128),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout127 (.I(net129),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout128 (.I(net129),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout129 (.I(net130),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout130 (.I(net131),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout131 (.I(net136),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout132 (.I(net134),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout133 (.I(net134),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout134 (.I(net135),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout135 (.I(net136),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout136 (.I(net137),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout137 (.I(net217),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout138 (.I(net141),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout139 (.I(net141),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout140 (.I(net141),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout141 (.I(net146),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout142 (.I(net144),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout143 (.I(net144),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout144 (.I(net146),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout145 (.I(net146),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout146 (.I(net153),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout147 (.I(net148),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout148 (.I(net152),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout149 (.I(net151),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout150 (.I(net151),
    .Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout151 (.I(net152),
    .Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout152 (.I(net153),
    .Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout153 (.I(net154),
    .Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout154 (.I(net178),
    .Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout155 (.I(net159),
    .Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout156 (.I(net157),
    .Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout157 (.I(net159),
    .Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout158 (.I(net177),
    .Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout159 (.I(net177),
    .Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout160 (.I(net161),
    .Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout161 (.I(net165),
    .Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout162 (.I(net165),
    .Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout163 (.I(net164),
    .Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout164 (.I(net165),
    .Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout165 (.I(net176),
    .Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout166 (.I(net169),
    .Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout167 (.I(net169),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout168 (.I(net169),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout169 (.I(net175),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout170 (.I(net171),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout171 (.I(net174),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout172 (.I(net173),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout173 (.I(net174),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout174 (.I(net175),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout175 (.I(net176),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout176 (.I(net177),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout177 (.I(net178),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout178 (.I(net216),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout179 (.I(net181),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout180 (.I(net181),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout181 (.I(net183),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout182 (.I(net183),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout183 (.I(net215),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout184 (.I(net186),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout185 (.I(net186),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout186 (.I(net189),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout187 (.I(net189),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout188 (.I(net189),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout189 (.I(net200),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout190 (.I(net194),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout191 (.I(net194),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout192 (.I(net194),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout193 (.I(net194),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout194 (.I(net199),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout195 (.I(net196),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout196 (.I(net198),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout197 (.I(net198),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout198 (.I(net199),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout199 (.I(net200),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout200 (.I(net214),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout201 (.I(net202),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout202 (.I(net204),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout203 (.I(net204),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout204 (.I(net213),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout205 (.I(net208),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout206 (.I(net208),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout207 (.I(net212),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout208 (.I(net212),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout209 (.I(net211),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout210 (.I(net211),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout211 (.I(net212),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout212 (.I(net213),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout213 (.I(net214),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout214 (.I(net215),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout215 (.I(net216),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout216 (.I(net217),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout217 (.I(net393),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout218 (.I(net220),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout219 (.I(net220),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout220 (.I(net222),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout221 (.I(net222),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout222 (.I(net228),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout223 (.I(net225),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout224 (.I(net225),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout225 (.I(net227),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout226 (.I(net227),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout227 (.I(net228),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout228 (.I(net234),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout229 (.I(net231),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout230 (.I(net231),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout231 (.I(net232),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout232 (.I(net234),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout233 (.I(net234),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout234 (.I(net241),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout235 (.I(net239),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout236 (.I(net239),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout237 (.I(net239),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout238 (.I(net239),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout239 (.I(net240),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout240 (.I(net241),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout241 (.I(net260),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout242 (.I(net243),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout243 (.I(net244),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout244 (.I(net250),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout245 (.I(net249),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout246 (.I(net249),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout247 (.I(net248),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout248 (.I(net249),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout249 (.I(net250),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout250 (.I(net258),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout251 (.I(net253),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout252 (.I(net253),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout253 (.I(net257),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout254 (.I(net255),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout255 (.I(net257),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout256 (.I(net257),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout257 (.I(net258),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout258 (.I(net259),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout259 (.I(net260),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout260 (.I(net286),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout261 (.I(net262),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout262 (.I(net285),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout263 (.I(net285),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout264 (.I(net267),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout265 (.I(net267),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout266 (.I(net267),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout267 (.I(net272),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout268 (.I(net271),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout269 (.I(net271),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout270 (.I(net271),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout271 (.I(net272),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout272 (.I(net273),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout273 (.I(net283),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout274 (.I(net276),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout275 (.I(net281),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout276 (.I(net281),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout277 (.I(net280),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout278 (.I(net280),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout279 (.I(net280),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout280 (.I(net281),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout281 (.I(net282),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout282 (.I(net283),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout283 (.I(net284),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout284 (.I(net285),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout285 (.I(net286),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout286 (.I(net392),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout287 (.I(net289),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout288 (.I(net290),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout289 (.I(net290),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout290 (.I(net295),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout291 (.I(net294),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout292 (.I(net294),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout293 (.I(net294),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout294 (.I(net295),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout295 (.I(net326),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout296 (.I(net300),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout297 (.I(net299),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout298 (.I(net299),
    .Z(net298));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout299 (.I(net300),
    .Z(net299));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout300 (.I(net310),
    .Z(net300));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout301 (.I(net304),
    .Z(net301));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout302 (.I(net304),
    .Z(net302));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout303 (.I(net304),
    .Z(net303));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout304 (.I(net309),
    .Z(net304));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout305 (.I(net307),
    .Z(net305));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout306 (.I(net307),
    .Z(net306));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout307 (.I(net308),
    .Z(net307));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout308 (.I(net309),
    .Z(net308));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout309 (.I(net310),
    .Z(net309));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout310 (.I(net325),
    .Z(net310));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout311 (.I(net312),
    .Z(net311));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout312 (.I(net319),
    .Z(net312));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout313 (.I(net319),
    .Z(net313));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout314 (.I(net318),
    .Z(net314));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout315 (.I(net318),
    .Z(net315));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout316 (.I(net318),
    .Z(net316));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout317 (.I(net318),
    .Z(net317));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout318 (.I(net319),
    .Z(net318));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout319 (.I(net324),
    .Z(net319));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout320 (.I(net322),
    .Z(net320));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout321 (.I(net322),
    .Z(net321));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout322 (.I(net324),
    .Z(net322));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout323 (.I(net324),
    .Z(net323));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout324 (.I(net325),
    .Z(net324));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout325 (.I(net326),
    .Z(net325));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout326 (.I(net391),
    .Z(net326));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout327 (.I(net328),
    .Z(net327));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout328 (.I(net329),
    .Z(net328));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout329 (.I(net333),
    .Z(net329));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout330 (.I(net333),
    .Z(net330));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout331 (.I(net332),
    .Z(net331));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout332 (.I(net333),
    .Z(net332));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout333 (.I(net338),
    .Z(net333));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout334 (.I(net336),
    .Z(net334));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout335 (.I(net336),
    .Z(net335));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout336 (.I(net337),
    .Z(net336));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout337 (.I(net338),
    .Z(net337));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout338 (.I(net353),
    .Z(net338));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout339 (.I(net343),
    .Z(net339));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout340 (.I(net343),
    .Z(net340));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout341 (.I(net343),
    .Z(net341));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout342 (.I(net343),
    .Z(net342));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout343 (.I(net352),
    .Z(net343));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout344 (.I(net347),
    .Z(net344));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout345 (.I(net347),
    .Z(net345));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout346 (.I(net347),
    .Z(net346));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout347 (.I(net351),
    .Z(net347));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout348 (.I(net350),
    .Z(net348));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout349 (.I(net351),
    .Z(net349));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout350 (.I(net351),
    .Z(net350));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout351 (.I(net352),
    .Z(net351));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout352 (.I(net353),
    .Z(net352));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout353 (.I(net367),
    .Z(net353));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout354 (.I(net356),
    .Z(net354));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout355 (.I(net360),
    .Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout356 (.I(net360),
    .Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout357 (.I(net359),
    .Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout358 (.I(net359),
    .Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout359 (.I(net360),
    .Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout360 (.I(net366),
    .Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout361 (.I(net364),
    .Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout362 (.I(net364),
    .Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout363 (.I(net365),
    .Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout364 (.I(net365),
    .Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout365 (.I(net366),
    .Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout366 (.I(net367),
    .Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout367 (.I(net390),
    .Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout368 (.I(net369),
    .Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout369 (.I(net374),
    .Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout370 (.I(net374),
    .Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout371 (.I(net373),
    .Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout372 (.I(net373),
    .Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout373 (.I(net374),
    .Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout374 (.I(net381),
    .Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout375 (.I(net376),
    .Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout376 (.I(net380),
    .Z(net376));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout377 (.I(net378),
    .Z(net377));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout378 (.I(net380),
    .Z(net378));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout379 (.I(net380),
    .Z(net379));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout380 (.I(net381),
    .Z(net380));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout381 (.I(net389),
    .Z(net381));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout382 (.I(net385),
    .Z(net382));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout383 (.I(net384),
    .Z(net383));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout384 (.I(net385),
    .Z(net384));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout385 (.I(net388),
    .Z(net385));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout386 (.I(net388),
    .Z(net386));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout387 (.I(net388),
    .Z(net387));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout388 (.I(net389),
    .Z(net388));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout389 (.I(net390),
    .Z(net389));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout390 (.I(net391),
    .Z(net390));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout391 (.I(net392),
    .Z(net391));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout392 (.I(net393),
    .Z(net392));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout393 (.I(net1),
    .Z(net393));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_394 (.ZN(net394));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__D (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__D (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__D (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__D (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A2 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__D (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__D (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A1 (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__D (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8528__D (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__D (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__D (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__D (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__D (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__D (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__D (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__D (.I(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__D (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__D (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8544__D (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__D (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__D (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__D (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__D (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__D (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__D (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__D (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__D (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__D (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__D (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__D (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__D (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__D (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__D (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__D (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__D (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__D (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__D (.I(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__D (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__D (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__D (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__D (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__B (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__I (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__I (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__I (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__I0 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__C (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__C (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__I (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__I (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__I (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__I0 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A3 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3969__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__I (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__B (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__B (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__I (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__I (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__B (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A1 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__I (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__I (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A3 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__B (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__I (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A3 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A3 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A3 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A3 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A3 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__B1 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__I0 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__I0 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__B1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__A3 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__I0 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__B1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__I (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__I1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__B2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__I0 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__I (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__S (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__S (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__S (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__B1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__S (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__S (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__I (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__B1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__B2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A3 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__I (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__S (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__S (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__S (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__S (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A3 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__B2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__I1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__B1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__C1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__B1 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__I (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__B2 (.I(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__B2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__B1 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__S (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4095__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__S (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__I0 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__I (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__C (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__C (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__I0 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__I (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A1 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__B2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__B1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__B1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__B1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__I (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__I (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__B1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A3 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__I (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__B (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A3 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A3 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A3 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__A2 (.I(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A2 (.I(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__B (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__A2 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__A2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A3 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A3 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A3 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A3 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A3 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4214__A2 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4176__A3 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A2 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A2 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__B2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__B (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A2 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A3 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__B (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__B1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__I0 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__B2 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A3 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__B1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A2 (.I(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__B2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A3 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A1 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A1 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__B (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__C (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A2 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A3 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A3 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A3 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__C (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__I (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A1 (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A3 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__B2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__B2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__B2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__I (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A2 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A4 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__I1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A3 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__B (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A4 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A4 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__C (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__C (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A2 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__B (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A3 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A3 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__I (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A3 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__B1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__B1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__B (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__C (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__A2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A2 (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A3 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A3 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A3 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__I (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A1 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A2 (.I(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__B1 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A4 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A3 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A2 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__A2 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A3 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A3 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__B1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A4 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__B2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A3 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__B (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A1 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__C (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__I (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__B (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__C (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A3 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__A1 (.I(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A3 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__I (.I(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A3 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__I (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A3 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A1 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__A1 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__B1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__B2 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A3 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__B2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__B (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A3 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A3 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__B2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__I (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A4 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__B (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A3 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__B1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__B (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__B (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__S (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A3 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A3 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__I0 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A1 (.I(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A2 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A2 (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__B (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A2 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A2 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__B2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A2 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A1 (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A2 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A2 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__C (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A3 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__B (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A3 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A2 (.I(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A3 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__S0 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__S0 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__I (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__I (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__C (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__I (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__B2 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A2 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__C (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__C (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__C (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__I (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__I (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__I (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__C (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__B (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__C (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__I (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__I (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__I (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__I (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__I (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__I (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__S (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__S (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__S (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__S (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__S (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__I2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__I (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__S (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__S (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__S (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__S (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__B1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__I3 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__I (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__I (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__I (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__A1 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__I (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__I (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__S0 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__S0 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__S0 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__I (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__S1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__S1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__S1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__S1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__B (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A2 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__I (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__B (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__B (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A2 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__I (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__I (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__I (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__I (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__I (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__I (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__S1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__S1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__B1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__I (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__I (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__I (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__S (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__I (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__S (.I(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__I (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A2 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__I (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__I (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__I (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__S (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__I (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__I (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__I (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__I (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__I (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__I (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__I (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__C (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__C (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A1 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__B2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__I (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__C (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__I (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__C (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__B (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__B (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__B2 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__I (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__I (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__I (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__I (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A1 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__I (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__S (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__I (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__S (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__S (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__S (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__I (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__I (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__I (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__I (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__B1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__S (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__S (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__S (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__S1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__S1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A1 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__B (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__I (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A2 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__I (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__I (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__I (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__I (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__I (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__I (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__S (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__B (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__I (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__I (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__I (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__I (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__I (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__I (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__I (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__I (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__I (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__B1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__S (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__S (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A2 (.I(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__I (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__I (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__I (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__I (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__I (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__S (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__S (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__S (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__B2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__B1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__S (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__S (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__B (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__B (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__C (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__B (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__C (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__C (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__C (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__I (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__I (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__B (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__C (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__B (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__B (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__B1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__I (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__C (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__C (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__C (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__B2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__I (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__B (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__C (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__B2 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__I0 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__I1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__B1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__B (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__B1 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__S (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__S (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__S (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__B1 (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__I (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__I (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__I (.I(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__S1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__S1 (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__C (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__B (.I(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__S (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__I (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__S (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__I (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__S (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__A2 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__I (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__I (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__C (.I(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__S (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__S (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__I (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__I (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A1 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A1 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A1 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__S1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__B (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__B (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__B (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__S1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__S1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__S1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__B (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A2 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A1 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__B (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__B (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__I (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__I (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__I (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__I (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__I (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__I (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__C (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__C (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__C (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__I (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__B (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__C (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__I (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__I (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__I (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__I (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A2 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__B (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__I (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__S (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__S (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A2 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__I0 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A1 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A2 (.I(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__I1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A2 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A2 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__I (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__I (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__I (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__I (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__I (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__I (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__I (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__S (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A1 (.I(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__S0 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__S0 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__I (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__S0 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__C (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__I (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__I (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__S (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__I0 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__I (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__I (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__I (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__S (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__B1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__I1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__S (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__I (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__I (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__S (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__I (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__I (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__I (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__S (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__S (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__S0 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__S (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__S (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__S (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__B2 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__B1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__B (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__C (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__I (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__I (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__B (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__B (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__I (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__B (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A1 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A2 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A2 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A1 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A1 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A1 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A2 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A2 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__S (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__S (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__S (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__I (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__S (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__B1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__B1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__B1 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A2 (.I(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__I0 (.I(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__I (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__S1 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__S1 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__I (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__B (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__B (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A1 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__B2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__I (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__S (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__S (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A2 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I0 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__B1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A1 (.I(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__S0 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__S (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A1 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__S (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A2 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__B (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__B (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__I (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I0 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__S (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__S (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__S (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__I (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__S (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__S1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A2 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I1 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__I (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__A1 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A2 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A2 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I2 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__S0 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__S (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I3 (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A2 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__C (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__S (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__I (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__I (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__B (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__B (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__B (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A1 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A1 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__S (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__S (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__S (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__B1 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__B1 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__B1 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__B2 (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__B2 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__B2 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__B2 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__S0 (.I(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A1 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A1 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A1 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__S (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__S (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__S (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__S (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__C (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__C (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__C (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__B (.I(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__I (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__I (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__S (.I(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__S (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__S (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A1 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__B (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__S (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__I (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__I (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A1 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A2 (.I(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A2 (.I(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__B (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__B (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__B (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__I (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__C (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__C (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__B (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__B (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__B (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__I1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__I3 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__I (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__I (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__I (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__S (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__S (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__S (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__S (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A2 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I0 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__S (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__S (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__S (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__S (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A2 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__S (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__S (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__S (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__S (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A2 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I2 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__I (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__S (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__S (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__S (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A2 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I3 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A1 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__S0 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__S0 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__S0 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__B (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A2 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__S (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__S (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__I (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__S (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__S (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__S (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__S (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__I0 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__I0 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__S (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__S (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__S (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__S (.I(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__S (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__S0 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__S0 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__S0 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A2 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__C (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__C (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A1 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__C (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__C (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__C (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__I1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__I3 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__I1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__I (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__S (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__S (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__S (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__S (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__S (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__S (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__I1 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__S (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__S (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__S (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__I2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__I3 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A1 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__S0 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__S0 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__S0 (.I(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__S (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__S0 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__S0 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__S0 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__I (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__I (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__I (.I(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__B2 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__S1 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__S1 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__S1 (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__S (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A2 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A2 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__S0 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__I1 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__B (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__B2 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__B2 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__B2 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__I (.I(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A1 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__B2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__S (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A2 (.I(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__B2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__I (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__I (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__S (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__I0 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__I1 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A2 (.I(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A3 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__I0 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A2 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__I1 (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__S (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__B2 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A1 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A1 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A2 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__A2 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__S (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__I (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__I (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A2 (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__I2 (.I(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A2 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__I3 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A2 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I1 (.I(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A1 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__S (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__S (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__S (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__S (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I3 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A2 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__I0 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__I0 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__I1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__I3 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I1 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__I3 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__I0 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__I0 (.I(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__I0 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__I3 (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A2 (.I(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A2 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I0 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__I3 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__I1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A2 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__B (.I(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__I (.I(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A2 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I0 (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A2 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I1 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I3 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A2 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__I0 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I0 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__I1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__I0 (.I(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I2 (.I(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__I0 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A2 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__I1 (.I(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A2 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__I3 (.I(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A2 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A2 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__I1 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__B (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__I (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__I (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__I (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__I (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__I (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__I (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__I (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__I (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__I (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A2 (.I(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A1 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__I (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__I (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__I (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A1 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__I (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__B2 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__I (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A1 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A1 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__I (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A1 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__B (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__I (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A2 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A2 (.I(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__B (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__I (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A2 (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__I (.I(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A3 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A3 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__I (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A3 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__C (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__C (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__C (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__I (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__S (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A1 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__I (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__I (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__S0 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__S0 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__I (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__I (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__B (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__C (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__C (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__I (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__I (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__I (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A2 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__B2 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__I (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__I (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__I (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__B2 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A1 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__I (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__C (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__B2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A3 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__B2 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A1 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A1 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A1 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A2 (.I(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__I (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__B (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__I (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A1 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__I (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__I (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__I (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__B (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__B (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__B (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__B2 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__C (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A2 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__S1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__S1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__I (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__I (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__I (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__C (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__I (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__C (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__C (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__I (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__B (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__I (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__I (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__B2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__I (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A2 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A2 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__B1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__B2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A2 (.I(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__B1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A2 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A2 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A1 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A2 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A2 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__B1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__I (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A2 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__B2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__B2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__B2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__B2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A2 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__B1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A2 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__I (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__I (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A3 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A3 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A2 (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A2 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A2 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__B1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A2 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__B1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__B1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__B1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__B1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__I (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__B1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__B2 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__I (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__I (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__B2 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__B1 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__B2 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__B2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__B2 (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__B2 (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__I (.I(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__S0 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__S0 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__S0 (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__C (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__C2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__C2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__B2 (.I(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__I (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__B2 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__I (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__B1 (.I(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__S (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__S (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__I (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__C (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A1 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A1 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A1 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A2 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__B2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A2 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__B1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__B1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__B1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__B1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__I (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__B (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__B1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__B1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__B1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__I (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__B2 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A1 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__C (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A1 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__I (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__B2 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__B2 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__B1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A2 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__A1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A1 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__I (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A1 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A1 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A1 (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__B (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__I (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__B (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A2 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A3 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A2 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__B2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__B2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__B2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__B2 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__C (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__S (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__I (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__I (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__B2 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__B2 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__B2 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__C (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__C (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__C (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__C (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__C (.I(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__C (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__C (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__C (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__S (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__B2 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__B2 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__B2 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__I (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__B (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__B (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__B (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__B (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__C (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__C (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__C (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6470__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A1 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__C (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__B (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__B (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__B (.I(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__S0 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A2 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A3 (.I(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__I (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__I (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__S (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A1 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__S0 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__B2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__A1 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A1 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__B2 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A1 (.I(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__B2 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__B (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__B (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__B (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A2 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A2 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A1 (.I(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A2 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A2 (.I(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__S (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__S (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__S (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A1 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__B2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__B2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__B2 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__S1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__A1 (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A2 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__B1 (.I(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__S (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A2 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__B1 (.I(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__I (.I(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A2 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__B1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__S (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__S (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__S (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__I (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__S1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A2 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__B1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__I (.I(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__I (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__I (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__B (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__B (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__I (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__I (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__B2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__B2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__I (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__I (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__B1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__C2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__B1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__B1 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__I (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__S (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__S (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__S (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__S (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__C1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__C1 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__C (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__C2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__C2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A2 (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__B1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__B1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__I (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__B1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__B2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__B2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A1 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__C2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__I (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__I (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__C (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__C (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A3 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__I (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__I (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__I (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__C (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A2 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__I (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__B (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__I (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__I (.I(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__B (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__B (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__S1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__S1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__S (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__S (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__B1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__B (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__I (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__I (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__I (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__I (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__B1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__B2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__B1 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__B2 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A2 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__I (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__I (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__I (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__B2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__B2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__B2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__C1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__B (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__B (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__I (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__I (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__S (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__B2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__B1 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__I (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A1 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__B2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A1 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__I (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__I (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A1 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A1 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__I (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__I (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__B (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__B (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__S (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__S (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A1 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__C (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__B (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__B (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A1 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__B2 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__B2 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__S (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__S (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__S (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A1 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__B2 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__B2 (.I(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A1 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__I (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__I (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__S (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A1 (.I(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__C (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__S1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__C (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A2 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A2 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__B1 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__B2 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__C1 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A2 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__C2 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A2 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__C2 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A2 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__B2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__C1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__C1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__B2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A1 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__B2 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__B2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__C1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__B1 (.I(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__C (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A1 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A1 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__B (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__B1 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__C (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__B2 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__C1 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__B2 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__C1 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__C1 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__C2 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__C2 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__C2 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__B2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__I (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__I (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__I (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__I (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__B1 (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__B1 (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A1 (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A2 (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__S (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__S (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__S (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__S (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__C1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__B1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__B2 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__B2 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__B (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__C (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__I (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__B2 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__I (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__I (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__C2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__C2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__S1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A1 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__B1 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__B2 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A1 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__C (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__B2 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__C (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__C (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A2 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__B2 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__B1 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__B1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__C1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__S (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__S (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__S (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__S (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__C1 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__C1 (.I(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A2 (.I(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A1 (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__B (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__B1 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__B1 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__B2 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__B1 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__B2 (.I(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__B2 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__C1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__B2 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__B1 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__B1 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__C (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__B2 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A2 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__B (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__I (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__B2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__B2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__C (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__C1 (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__B2 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__B1 (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__C2 (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__C2 (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__B (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A3 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A4 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A3 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__B1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__B2 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A2 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A1 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A1 (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A1 (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__S (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__S (.I(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__C1 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A2 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A1 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A1 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A1 (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__S (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__S (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__B1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__B1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A2 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A1 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__I (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__B1 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__B1 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__B2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__B2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__C1 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__B1 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__B1 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__B1 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__B2 (.I(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__B2 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A2 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__C1 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__B1 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__A2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__B1 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__C (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__I (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A1 (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__I (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__B2 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A2 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__B1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A2 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__B (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A3 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A2 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A1 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__S0 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A1 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__B (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__B1 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__B1 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A4 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__A1 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A1 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__B2 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__C1 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__B2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__B1 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A2 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A2 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__B1 (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__B1 (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__C (.I(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__B1 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A2 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__B (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A3 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A2 (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A2 (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A3 (.I(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__B1 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A1 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A1 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__I (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__I (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A2 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A2 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A1 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A1 (.I(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A2 (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__I (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__I (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__I (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__I (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__C (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__I (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A1 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A2 (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__C (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__C (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__I (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__B (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__C (.I(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__I (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A2 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__I (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__B (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__B (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A1 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__I (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__I (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__I (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__I (.I(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A1 (.I(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A1 (.I(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__C (.I(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A2 (.I(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__S (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__I (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__I (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__I (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__I (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A1 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__I (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__I (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A3 (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A1 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A3 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A1 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__B (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__C (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__C (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__C (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__B1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__B1 (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__B (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__B (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A1 (.I(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__B (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__B (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__B (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__C (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6118__A2 (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__B2 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__B (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__C (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__C (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__C (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__B (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__S1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A2 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A2 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A2 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__B (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__B (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__C (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__C (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__A2 (.I(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A1 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__B (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A1 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__B2 (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__B (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__B (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__B (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__B (.I(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__S1 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__S1 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__S1 (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__C (.I(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A2 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__B (.I(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__B (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A1 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A1 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A2 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__B1 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__I (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__I (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__C (.I(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__C (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__C (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A1 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A1 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__B (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__B1 (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__B (.I(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__B1 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A1 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A1 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A1 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__B (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__B (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__B (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__B (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A1 (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A1 (.I(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A1 (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__I (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__I (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__B2 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A2 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__B1 (.I(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A1 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__B2 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__B2 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__B2 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A1 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A2 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__S (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__S (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__S (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__S (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__B2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__B2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__B2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__B2 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A2 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__A2 (.I(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A2 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A2 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A2 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__I3 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A2 (.I(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A2 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__C (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__I3 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A1 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__C (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__B1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__B2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__B1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__B1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__B1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__C2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__B2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__C2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__B2 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__B1 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__B1 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__C (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__C (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__C (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__C (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A1 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A1 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A1 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__B2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__B2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__I (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__B1 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__C2 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__C2 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__C2 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__B2 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__B1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__B1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__B1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__C1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__B1 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A1 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__B2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A1 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A1 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A1 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A3 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__B1 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A2 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__B2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__I (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__C2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__B (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__B2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__B1 (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A1 (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__C1 (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__B (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__B2 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__B2 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__B2 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__B1 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__B (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A3 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A1 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__B (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A1 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__B (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__C (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A2 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__B (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__B (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__B (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__B (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__B (.I(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A2 (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A3 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__B1 (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__A2 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A4 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A3 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__I (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__I (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__I (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__I (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__I0 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__I0 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__I0 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__I0 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A2 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A2 (.I(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__I (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__S (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__S (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__S (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__S (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__I0 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__I0 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__I0 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__I0 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__I (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__I0 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__I0 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__I0 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__I0 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__I0 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__I0 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__I0 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__I0 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__I0 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__I0 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__I0 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__I0 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__S (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__S (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__S (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__S (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__I (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__I0 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__I0 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__I0 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__I0 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__I0 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__I0 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__I0 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__I0 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__I0 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__I0 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__I0 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__I0 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A1 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A1 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A1 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__S (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__S (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__S (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__S (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__S (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__S (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__S (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__S (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__I (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__I (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__I (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__I (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__I0 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__I0 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__I1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__I1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A2 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__A3 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A2 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__I (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__I (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__S (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__S (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__S (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__S (.I(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__I (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__I0 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__I0 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__I1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__I1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__I (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7472__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__I0 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__I0 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__I0 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__I1 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__I (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__I0 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A1 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__I1 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__I1 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__I1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__I1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__I0 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__I1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__I1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__I0 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__I1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__I1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A3 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A3 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A3 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__S (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__I (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__I (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A2 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__S (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__S (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__S (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A3 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__I (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6902__I (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__I0 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__I0 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__I0 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__I0 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__A3 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__A3 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A3 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A3 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__I (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__I (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__S (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__S (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__S (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__S (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__I0 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__I0 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__I0 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__I0 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__I0 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__I0 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__I0 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__I0 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__I0 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__I0 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__I0 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__I0 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__S (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__S (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__S (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__S (.I(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__I0 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__I0 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__I0 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I0 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__I0 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__I0 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__I0 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__I0 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__A1 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A3 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__I (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__I (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__S (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__S (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__S (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__S (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__S (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__S (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__S (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__S (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__I0 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__I0 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__I0 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__I0 (.I(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__I (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__I (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__S (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__S (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__S (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__S (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__S (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__S (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__S (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6983__S (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__I (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__I (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__S (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__S (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__S (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__S (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__S (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__S (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__S (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__S (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__I0 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__I0 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__I0 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__I0 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A3 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A3 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__I (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__I (.I(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__S (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__S (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__S (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__S (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__I0 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__I0 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__I0 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__I0 (.I(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__I0 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__I0 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__I0 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__I0 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__I0 (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__I0 (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__I0 (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__I0 (.I(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__I0 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__I0 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__I0 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__I0 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__S (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__S (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__S (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__S (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__I0 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__I0 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__I0 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__I0 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__I0 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__I0 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__I0 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__I0 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__S (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A2 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A2 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__S (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__S (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__S (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__S (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__S (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__S (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__I (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__I (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__S (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__S (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__S (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__S (.I(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__S (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__S (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__S (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__S (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__I0 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__I0 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__I0 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__I0 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__I (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__I (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__S (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__S (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__S (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__S (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__I0 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__I0 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__I0 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__I0 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__I (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__I (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__S (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__S (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__S (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__S (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__I0 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__I0 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__I0 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__I0 (.I(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I0 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__I0 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__I0 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__I0 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__I0 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__I0 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__I0 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__I0 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__I0 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I0 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__I0 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__I0 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__S (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__S (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__S (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__S (.I(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__I0 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__I0 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__I0 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I0 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__I0 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__I0 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__I0 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__I0 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__S (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__I (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__I (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__S (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__S (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__S (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__S (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__I1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__I (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__I (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__S (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__S (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__S (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__S (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__S (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__S (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__S (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__S (.I(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__I0 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__I0 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__I0 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__I0 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__I (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__I (.I(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__S (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__S (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__S (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__S (.I(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__I (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__I (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__S (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__S (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__S (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__S (.I(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__S (.I(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__I0 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__I0 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__I0 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__I0 (.I(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__I (.I(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__I (.I(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__S (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A2 (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__S (.I(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__S (.I(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__S (.I(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__S (.I(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__I (.I(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__A2 (.I(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A1 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A1 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A1 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__A1 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A1 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A1 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A1 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A1 (.I(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__I0 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__I0 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__I0 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__I0 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__I0 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__I0 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__I0 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__I0 (.I(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__I0 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__I0 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__I0 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__I0 (.I(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__I (.I(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__S (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A2 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A2 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__S (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__S (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__S (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__S (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__I (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A2 (.I(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__I (.I(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__S (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__S (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__S (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__S (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__I0 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__I0 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__I0 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__I0 (.I(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__S (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__S (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__S (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__S (.I(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__I0 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__I0 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__I0 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__I0 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__I (.I(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__I (.I(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__S (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__S (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__S (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__S (.I(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__I0 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__I0 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__I0 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__I0 (.I(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__I0 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__I0 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__I0 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__I0 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__I (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__I (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__S (.I(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__S (.I(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__S (.I(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__S (.I(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__I0 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__I0 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__I0 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__I0 (.I(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__S (.I(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__I0 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__I0 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__I0 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__I0 (.I(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__I0 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__I0 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__I0 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__I0 (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__I (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__I (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__S (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__S (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__S (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__S (.I(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__S (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__S (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__S (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__S (.I(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__I (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__I (.I(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__S (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__S (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__S (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__S (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__I0 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__I0 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__I0 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__I0 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__I0 (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__I0 (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__I0 (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__I0 (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__S (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__S (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__S (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__S (.I(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__I0 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__I0 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__I0 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__I0 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__S (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__S (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__I (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__I (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__S (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__S (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__S (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__S (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7555__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__A2 (.I(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__I0 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__I0 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__I0 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__I0 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__I0 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__I0 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__I0 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__I0 (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__I (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__I (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__S (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__S (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__S (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__S (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__I0 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__I0 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__I0 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__I0 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__S (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__S (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__S (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__S (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__I0 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__I0 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__I0 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__I0 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__I0 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__I0 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__I0 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__I0 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__S (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__S (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__I (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__I (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__S (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__S (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__S (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__S (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7600__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__I (.I(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__I (.I(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A2 (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__A2 (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__S (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__S (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__S (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__I (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__S (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__S (.I(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__A2 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A2 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A2 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A2 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__I0 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__I0 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__I0 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__I0 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__I (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__I (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__S (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__S (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__S (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__S (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__I (.I(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__I (.I(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__S (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__S (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__S (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__S (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__I (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__I (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__I (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__I (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__S (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__S (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__S (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__S (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__I (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__S (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__S (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__S (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__S (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A1 (.I(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A1 (.I(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A1 (.I(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A1 (.I(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__I (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__I (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__A2 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A2 (.I(\mod.Arithmetic.ACTI.x[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__I (.I(\mod.Arithmetic.ACTI.x[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__B (.I(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__A2 (.I(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__I (.I(\mod.Arithmetic.ACTI.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__C (.I(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A2 (.I(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__I (.I(\mod.Arithmetic.ACTI.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A2 (.I(\mod.Arithmetic.ACTI.x[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A2 (.I(\mod.Arithmetic.ACTI.x[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__I (.I(\mod.Arithmetic.ACTI.x[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__C (.I(\mod.Arithmetic.ACTI.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__A2 (.I(\mod.Arithmetic.ACTI.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__I (.I(\mod.Arithmetic.ACTI.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__C (.I(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A2 (.I(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__I (.I(\mod.Arithmetic.ACTI.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A2 (.I(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__B2 (.I(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__B2 (.I(\mod.Arithmetic.ACTI.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I0 (.I(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A2 (.I(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__I (.I(\mod.Arithmetic.ACTI.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__I (.I(\mod.Arithmetic.CN.F_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__I (.I(\mod.Arithmetic.CN.F_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__I (.I(\mod.Arithmetic.CN.F_in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__I (.I(\mod.Arithmetic.CN.I_in[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__I (.I(\mod.Arithmetic.CN.I_in[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A2 (.I(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__I0 (.I(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__I (.I(\mod.Arithmetic.CN.I_in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__I (.I(\mod.Arithmetic.CN.I_in[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__I (.I(\mod.Arithmetic.CN.I_in[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A2 (.I(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__I (.I(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__I (.I(\mod.Arithmetic.CN.I_in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__I (.I(\mod.Arithmetic.CN.I_in[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__I (.I(\mod.Arithmetic.CN.I_in[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(\mod.Arithmetic.CN.I_in[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A1 (.I(\mod.Arithmetic.CN.I_in[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__I (.I(\mod.Arithmetic.CN.I_in[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A2 (.I(\mod.Arithmetic.CN.I_in[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__I (.I(\mod.Arithmetic.CN.I_in[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(\mod.Arithmetic.CN.I_in[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__I0 (.I(\mod.Arithmetic.CN.I_in[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__I (.I(\mod.Arithmetic.CN.I_in[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A2 (.I(\mod.Arithmetic.CN.I_in[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__I (.I(\mod.Arithmetic.CN.I_in[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A3 (.I(\mod.Arithmetic.CN.I_in[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(\mod.Arithmetic.CN.I_in[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__I (.I(\mod.Arithmetic.CN.I_in[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A3 (.I(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A2 (.I(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A2 (.I(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__I (.I(\mod.Arithmetic.CN.I_in[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A2 (.I(\mod.Arithmetic.CN.I_in[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__I (.I(\mod.Arithmetic.CN.I_in[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(\mod.Arithmetic.CN.I_in[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__B2 (.I(\mod.Arithmetic.CN.I_in[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__I (.I(\mod.Arithmetic.CN.I_in[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A1 (.I(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__I (.I(\mod.Arithmetic.CN.I_in[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A2 (.I(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A2 (.I(\mod.Arithmetic.CN.I_in[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(\mod.Arithmetic.CN.I_in[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A2 (.I(\mod.Arithmetic.CN.I_in[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__I (.I(\mod.Arithmetic.CN.I_in[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A2 (.I(\mod.Arithmetic.CN.I_in[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__I (.I(\mod.Arithmetic.CN.I_in[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(\mod.Arithmetic.CN.I_in[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__I (.I(\mod.Arithmetic.CN.I_in[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__I (.I(\mod.Arithmetic.CN.I_in[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(\mod.Arithmetic.CN.I_in[32] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__B2 (.I(\mod.Arithmetic.CN.I_in[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A3 (.I(\mod.Arithmetic.CN.I_in[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A2 (.I(\mod.Arithmetic.CN.I_in[33] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__I (.I(\mod.Arithmetic.CN.I_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A2 (.I(\mod.Arithmetic.CN.I_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A1 (.I(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(\mod.Arithmetic.CN.I_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(\mod.Arithmetic.CN.I_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__I (.I(\mod.Arithmetic.CN.I_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__A1 (.I(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__I (.I(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(\mod.Arithmetic.CN.I_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(\mod.Arithmetic.CN.I_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(\mod.Arithmetic.CN.I_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(\mod.Arithmetic.CN.I_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(\mod.Arithmetic.CN.I_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A2 (.I(\mod.Arithmetic.CN.I_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__I (.I(\mod.Arithmetic.CN.I_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A2 (.I(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__B2 (.I(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__A3 (.I(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A2 (.I(\mod.Arithmetic.CN.I_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__I (.I(\mod.Arithmetic.CN.I_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(\mod.Arithmetic.CN.I_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(\mod.Arithmetic.CN.I_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A2 (.I(\mod.Arithmetic.CN.I_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(\mod.Arithmetic.CN.I_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__I (.I(\mod.Arithmetic.CN.I_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A2 (.I(\mod.Arithmetic.CN.I_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(\mod.Arithmetic.CN.I_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(\mod.Arithmetic.CN.I_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(\mod.Arithmetic.CN.I_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A2 (.I(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A2 (.I(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A1 (.I(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(\mod.Arithmetic.CN.I_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(\mod.Arithmetic.CN.I_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(\mod.Arithmetic.CN.I_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(\mod.Arithmetic.CN.I_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__I (.I(\mod.Arithmetic.CN.I_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(\mod.Arithmetic.CN.I_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(\mod.Arithmetic.CN.I_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A2 (.I(\mod.Arithmetic.CN.I_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__A3 (.I(\mod.Arithmetic.CN.I_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A1 (.I(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A1 (.I(\mod.Arithmetic.CN.I_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(\mod.Arithmetic.CN.I_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(\mod.Arithmetic.CN.I_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__A2 (.I(\mod.Arithmetic.CN.I_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A2 (.I(\mod.Arithmetic.CN.I_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A2 (.I(\mod.Arithmetic.CN.I_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__I (.I(\mod.Arithmetic.CN.I_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__A2 (.I(\mod.Arithmetic.CN.I_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__I (.I(\mod.Arithmetic.CN.I_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A3 (.I(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A1 (.I(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__I (.I(\mod.Arithmetic.CN.I_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A3 (.I(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A2 (.I(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A3 (.I(\mod.Arithmetic.CN.I_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(\mod.Arithmetic.CN.I_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A2 (.I(\mod.Arithmetic.CN.I_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(\mod.Arithmetic.CN.I_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A1 (.I(\mod.Arithmetic.CN.I_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A2 (.I(\mod.Arithmetic.CN.I_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(\mod.Arithmetic.CN.I_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(\mod.Arithmetic.CN.I_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A2 (.I(\mod.Arithmetic.CN.I_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(\mod.Arithmetic.CN.I_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A2 (.I(\mod.Arithmetic.CN.I_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A2 (.I(\mod.Arithmetic.CN.I_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A2 (.I(\mod.Arithmetic.CN.I_in[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__I1 (.I(\mod.Arithmetic.CN.I_in[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A2 (.I(\mod.Arithmetic.CN.I_in[70] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(\mod.Arithmetic.CN.I_in[71] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A1 (.I(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__A2 (.I(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__I (.I(\mod.Arithmetic.CN.I_in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A4 (.I(\mod.Arithmetic.CN.I_in[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__I (.I(\mod.Arithmetic.CN.I_in[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__I (.I(\mod.Arithmetic.I_out[72] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__I1 (.I(\mod.Arithmetic.I_out[72] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__B (.I(\mod.Arithmetic.I_out[72] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__I1 (.I(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__I (.I(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__B2 (.I(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(\mod.Arithmetic.I_out[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A3 (.I(\mod.Arithmetic.I_out[79] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A2 (.I(\mod.Arithmetic.I_out[79] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__I (.I(\mod.Arithmetic.I_out[79] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A2 (.I(\mod.Arithmetic.I_out[79] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__I0 (.I(\mod.Data_Mem.F_M.MRAM[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__B2 (.I(\mod.Data_Mem.F_M.MRAM[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__I0 (.I(\mod.Data_Mem.F_M.MRAM[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I2 (.I(\mod.Data_Mem.F_M.MRAM[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A2 (.I(\mod.Data_Mem.F_M.MRAM[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__I1 (.I(\mod.Data_Mem.F_M.MRAM[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(\mod.Data_Mem.F_M.MRAM[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__I0 (.I(\mod.Data_Mem.F_M.MRAM[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__I1 (.I(\mod.Data_Mem.F_M.MRAM[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A2 (.I(\mod.Data_Mem.F_M.MRAM[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__B2 (.I(\mod.Data_Mem.F_M.MRAM[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__I1 (.I(\mod.Data_Mem.F_M.MRAM[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A2 (.I(\mod.Data_Mem.F_M.MRAM[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(\mod.Data_Mem.F_M.MRAM[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__B1 (.I(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A2 (.I(\mod.Data_Mem.F_M.MRAM[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__B1 (.I(\mod.Data_Mem.F_M.MRAM[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__I1 (.I(\mod.Data_Mem.F_M.MRAM[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__B1 (.I(\mod.Data_Mem.F_M.MRAM[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__I0 (.I(\mod.Data_Mem.F_M.MRAM[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__B1 (.I(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(\mod.Data_Mem.F_M.MRAM[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__B1 (.I(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__B2 (.I(\mod.Data_Mem.F_M.MRAM[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__B1 (.I(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__B2 (.I(\mod.Data_Mem.F_M.MRAM[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__B1 (.I(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(\mod.Data_Mem.F_M.MRAM[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__A2 (.I(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(\mod.Data_Mem.F_M.MRAM[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A2 (.I(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A1 (.I(\mod.Data_Mem.F_M.MRAM[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A2 (.I(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__I1 (.I(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(\mod.Data_Mem.F_M.MRAM[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__I0 (.I(\mod.Data_Mem.F_M.MRAM[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__I1 (.I(\mod.Data_Mem.F_M.MRAM[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__I1 (.I(\mod.Data_Mem.F_M.MRAM[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__I0 (.I(\mod.Data_Mem.F_M.MRAM[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I0 (.I(\mod.Data_Mem.F_M.MRAM[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(\mod.Data_Mem.F_M.MRAM[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A2 (.I(\mod.Data_Mem.F_M.MRAM[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I1 (.I(\mod.Data_Mem.F_M.MRAM[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7132__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A2 (.I(\mod.Data_Mem.F_M.MRAM[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__I1 (.I(\mod.Data_Mem.F_M.MRAM[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A2 (.I(\mod.Data_Mem.F_M.MRAM[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I0 (.I(\mod.Data_Mem.F_M.MRAM[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(\mod.Data_Mem.F_M.MRAM[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__B2 (.I(\mod.Data_Mem.F_M.MRAM[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A2 (.I(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A2 (.I(\mod.Data_Mem.F_M.MRAM[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(\mod.Data_Mem.F_M.MRAM[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__I1 (.I(\mod.Data_Mem.F_M.MRAM[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(\mod.Data_Mem.F_M.MRAM[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__I0 (.I(\mod.Data_Mem.F_M.MRAM[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__I (.I(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A3 (.I(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__I2 (.I(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__I1 (.I(\mod.Data_Mem.F_M.MRAM[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__I (.I(\mod.Data_Mem.F_M.MRAM[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(\mod.Data_Mem.F_M.MRAM[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I1 (.I(\mod.Data_Mem.F_M.MRAM[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__I (.I(\mod.Data_Mem.F_M.MRAM[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A2 (.I(\mod.Data_Mem.F_M.MRAM[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__I1 (.I(\mod.Data_Mem.F_M.MRAM[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__I (.I(\mod.Data_Mem.F_M.MRAM[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(\mod.Data_Mem.F_M.MRAM[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__I1 (.I(\mod.Data_Mem.F_M.MRAM[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__I (.I(\mod.Data_Mem.F_M.MRAM[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A2 (.I(\mod.Data_Mem.F_M.MRAM[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__I1 (.I(\mod.Data_Mem.F_M.MRAM[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__I (.I(\mod.Data_Mem.F_M.MRAM[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__I3 (.I(\mod.Data_Mem.F_M.MRAM[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__I0 (.I(\mod.Data_Mem.F_M.MRAM[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__I (.I(\mod.Data_Mem.F_M.MRAM[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__I3 (.I(\mod.Data_Mem.F_M.MRAM[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__I0 (.I(\mod.Data_Mem.F_M.MRAM[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__I (.I(\mod.Data_Mem.F_M.MRAM[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A2 (.I(\mod.Data_Mem.F_M.MRAM[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I0 (.I(\mod.Data_Mem.F_M.MRAM[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__I (.I(\mod.Data_Mem.F_M.MRAM[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A2 (.I(\mod.Data_Mem.F_M.MRAM[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__I0 (.I(\mod.Data_Mem.F_M.MRAM[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__I (.I(\mod.Data_Mem.F_M.MRAM[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A2 (.I(\mod.Data_Mem.F_M.MRAM[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__I0 (.I(\mod.Data_Mem.F_M.MRAM[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__I (.I(\mod.Data_Mem.F_M.MRAM[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(\mod.Data_Mem.F_M.MRAM[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__I0 (.I(\mod.Data_Mem.F_M.MRAM[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__I (.I(\mod.Data_Mem.F_M.MRAM[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(\mod.Data_Mem.F_M.MRAM[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A1 (.I(\mod.Data_Mem.F_M.MRAM[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__I (.I(\mod.Data_Mem.F_M.MRAM[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__A1 (.I(\mod.Data_Mem.F_M.MRAM[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__I (.I(\mod.Data_Mem.F_M.MRAM[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__B1 (.I(\mod.Data_Mem.F_M.MRAM[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__I1 (.I(\mod.Data_Mem.F_M.MRAM[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A2 (.I(\mod.Data_Mem.F_M.MRAM[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__B2 (.I(\mod.Data_Mem.F_M.MRAM[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__I1 (.I(\mod.Data_Mem.F_M.MRAM[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A2 (.I(\mod.Data_Mem.F_M.MRAM[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A1 (.I(\mod.Data_Mem.F_M.MRAM[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A2 (.I(\mod.Data_Mem.F_M.MRAM[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I3 (.I(\mod.Data_Mem.F_M.MRAM[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A2 (.I(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A2 (.I(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__I0 (.I(\mod.Data_Mem.F_M.MRAM[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__I1 (.I(\mod.Data_Mem.F_M.MRAM[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__I0 (.I(\mod.Data_Mem.F_M.MRAM[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__I0 (.I(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__I0 (.I(\mod.Data_Mem.F_M.MRAM[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I0 (.I(\mod.Data_Mem.F_M.MRAM[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__B1 (.I(\mod.Data_Mem.F_M.MRAM[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__B1 (.I(\mod.Data_Mem.F_M.MRAM[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__B1 (.I(\mod.Data_Mem.F_M.MRAM[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__I1 (.I(\mod.Data_Mem.F_M.MRAM[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__B1 (.I(\mod.Data_Mem.F_M.MRAM[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A2 (.I(\mod.Data_Mem.F_M.MRAM[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__B1 (.I(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__I1 (.I(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__B1 (.I(\mod.Data_Mem.F_M.MRAM[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I (.I(\mod.Data_Mem.F_M.MRAM[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__B1 (.I(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__I1 (.I(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I1 (.I(\mod.Data_Mem.F_M.MRAM[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__B1 (.I(\mod.Data_Mem.F_M.MRAM[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A1 (.I(\mod.Data_Mem.F_M.MRAM[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(\mod.Data_Mem.F_M.MRAM[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A1 (.I(\mod.Data_Mem.F_M.MRAM[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__I0 (.I(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A2 (.I(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(\mod.Data_Mem.F_M.MRAM[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A2 (.I(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(\mod.Data_Mem.F_M.MRAM[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I2 (.I(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A2 (.I(\mod.Data_Mem.F_M.MRAM[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__I1 (.I(\mod.Data_Mem.F_M.MRAM[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__I0 (.I(\mod.Data_Mem.F_M.MRAM[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__I (.I(\mod.Data_Mem.F_M.MRAM[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__I0 (.I(\mod.Data_Mem.F_M.MRAM[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__I (.I(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I3 (.I(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__I0 (.I(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__I (.I(\mod.Data_Mem.F_M.MRAM[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A2 (.I(\mod.Data_Mem.F_M.MRAM[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__I (.I(\mod.Data_Mem.F_M.MRAM[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A2 (.I(\mod.Data_Mem.F_M.MRAM[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__I1 (.I(\mod.Data_Mem.F_M.MRAM[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__I (.I(\mod.Data_Mem.F_M.MRAM[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__I1 (.I(\mod.Data_Mem.F_M.MRAM[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__I0 (.I(\mod.Data_Mem.F_M.MRAM[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__I (.I(\mod.Data_Mem.F_M.MRAM[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__I1 (.I(\mod.Data_Mem.F_M.MRAM[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I0 (.I(\mod.Data_Mem.F_M.MRAM[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__I (.I(\mod.Data_Mem.F_M.MRAM[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(\mod.Data_Mem.F_M.MRAM[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__I0 (.I(\mod.Data_Mem.F_M.MRAM[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__I (.I(\mod.Data_Mem.F_M.MRAM[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A2 (.I(\mod.Data_Mem.F_M.MRAM[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__I0 (.I(\mod.Data_Mem.F_M.MRAM[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__I (.I(\mod.Data_Mem.F_M.MRAM[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A2 (.I(\mod.Data_Mem.F_M.MRAM[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__I0 (.I(\mod.Data_Mem.F_M.MRAM[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__I (.I(\mod.Data_Mem.F_M.MRAM[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A2 (.I(\mod.Data_Mem.F_M.MRAM[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(\mod.Data_Mem.F_M.MRAM[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__I (.I(\mod.Data_Mem.F_M.MRAM[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(\mod.Data_Mem.F_M.MRAM[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A2 (.I(\mod.Data_Mem.F_M.MRAM[768][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I1 (.I(\mod.Data_Mem.F_M.MRAM[768][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__I0 (.I(\mod.Data_Mem.F_M.MRAM[769][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A2 (.I(\mod.Data_Mem.F_M.MRAM[769][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__I0 (.I(\mod.Data_Mem.F_M.MRAM[769][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__I1 (.I(\mod.Data_Mem.F_M.MRAM[769][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__B2 (.I(\mod.Data_Mem.F_M.MRAM[769][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I0 (.I(\mod.Data_Mem.F_M.MRAM[769][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__I0 (.I(\mod.Data_Mem.F_M.MRAM[770][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__I0 (.I(\mod.Data_Mem.F_M.MRAM[770][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__I0 (.I(\mod.Data_Mem.F_M.MRAM[770][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__I0 (.I(\mod.Data_Mem.F_M.MRAM[770][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I1 (.I(\mod.Data_Mem.F_M.MRAM[770][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__I0 (.I(\mod.Data_Mem.F_M.MRAM[771][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A2 (.I(\mod.Data_Mem.F_M.MRAM[771][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A2 (.I(\mod.Data_Mem.F_M.MRAM[771][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(\mod.Data_Mem.F_M.MRAM[771][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A2 (.I(\mod.Data_Mem.F_M.MRAM[771][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A2 (.I(\mod.Data_Mem.F_M.MRAM[771][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A2 (.I(\mod.Data_Mem.F_M.MRAM[771][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__I0 (.I(\mod.Data_Mem.F_M.MRAM[771][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I0 (.I(\mod.Data_Mem.F_M.MRAM[771][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__I0 (.I(\mod.Data_Mem.F_M.MRAM[771][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6032__I1 (.I(\mod.Data_Mem.F_M.MRAM[771][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I0 (.I(\mod.Data_Mem.F_M.MRAM[771][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__I (.I(\mod.Data_Mem.F_M.MRAM[772][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A2 (.I(\mod.Data_Mem.F_M.MRAM[772][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__I1 (.I(\mod.Data_Mem.F_M.MRAM[772][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__I (.I(\mod.Data_Mem.F_M.MRAM[772][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A2 (.I(\mod.Data_Mem.F_M.MRAM[772][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I1 (.I(\mod.Data_Mem.F_M.MRAM[772][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__I (.I(\mod.Data_Mem.F_M.MRAM[772][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A2 (.I(\mod.Data_Mem.F_M.MRAM[772][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__I1 (.I(\mod.Data_Mem.F_M.MRAM[772][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__I (.I(\mod.Data_Mem.F_M.MRAM[773][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(\mod.Data_Mem.F_M.MRAM[773][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__I0 (.I(\mod.Data_Mem.F_M.MRAM[773][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__I (.I(\mod.Data_Mem.F_M.MRAM[773][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A2 (.I(\mod.Data_Mem.F_M.MRAM[773][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__I0 (.I(\mod.Data_Mem.F_M.MRAM[773][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__I (.I(\mod.Data_Mem.F_M.MRAM[773][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A2 (.I(\mod.Data_Mem.F_M.MRAM[773][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__I0 (.I(\mod.Data_Mem.F_M.MRAM[773][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__I (.I(\mod.Data_Mem.F_M.MRAM[773][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A2 (.I(\mod.Data_Mem.F_M.MRAM[773][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__I0 (.I(\mod.Data_Mem.F_M.MRAM[773][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__I (.I(\mod.Data_Mem.F_M.MRAM[773][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A2 (.I(\mod.Data_Mem.F_M.MRAM[773][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__I0 (.I(\mod.Data_Mem.F_M.MRAM[773][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__I (.I(\mod.Data_Mem.F_M.MRAM[775][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(\mod.Data_Mem.F_M.MRAM[775][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A2 (.I(\mod.Data_Mem.F_M.MRAM[780][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A2 (.I(\mod.Data_Mem.F_M.MRAM[780][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__B2 (.I(\mod.Data_Mem.F_M.MRAM[780][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(\mod.Data_Mem.F_M.MRAM[780][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__B2 (.I(\mod.Data_Mem.F_M.MRAM[780][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A2 (.I(\mod.Data_Mem.F_M.MRAM[780][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__I0 (.I(\mod.Data_Mem.F_M.MRAM[780][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__B2 (.I(\mod.Data_Mem.F_M.MRAM[780][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A2 (.I(\mod.Data_Mem.F_M.MRAM[780][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__B2 (.I(\mod.Data_Mem.F_M.MRAM[780][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A2 (.I(\mod.Data_Mem.F_M.MRAM[780][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__B2 (.I(\mod.Data_Mem.F_M.MRAM[780][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7482__I1 (.I(\mod.Data_Mem.F_M.MRAM[780][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A1 (.I(\mod.Data_Mem.F_M.MRAM[780][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__B2 (.I(\mod.Data_Mem.F_M.MRAM[780][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A2 (.I(\mod.Data_Mem.F_M.MRAM[781][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A2 (.I(\mod.Data_Mem.F_M.MRAM[781][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A2 (.I(\mod.Data_Mem.F_M.MRAM[781][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A2 (.I(\mod.Data_Mem.F_M.MRAM[781][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__I (.I(\mod.Data_Mem.F_M.MRAM[781][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__I2 (.I(\mod.Data_Mem.F_M.MRAM[781][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A2 (.I(\mod.Data_Mem.F_M.MRAM[781][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__A2 (.I(\mod.Data_Mem.F_M.MRAM[781][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__I1 (.I(\mod.Data_Mem.F_M.MRAM[781][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A1 (.I(\mod.Data_Mem.F_M.MRAM[781][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A2 (.I(\mod.Data_Mem.F_M.MRAM[782][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__I0 (.I(\mod.Data_Mem.F_M.MRAM[782][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__B1 (.I(\mod.Data_Mem.F_M.MRAM[782][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__I0 (.I(\mod.Data_Mem.F_M.MRAM[782][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7513__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__B1 (.I(\mod.Data_Mem.F_M.MRAM[782][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__I0 (.I(\mod.Data_Mem.F_M.MRAM[782][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__B1 (.I(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__I0 (.I(\mod.Data_Mem.F_M.MRAM[782][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B1 (.I(\mod.Data_Mem.F_M.MRAM[782][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A2 (.I(\mod.Data_Mem.F_M.MRAM[782][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__B1 (.I(\mod.Data_Mem.F_M.MRAM[782][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A2 (.I(\mod.Data_Mem.F_M.MRAM[782][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__I1 (.I(\mod.Data_Mem.F_M.MRAM[782][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__B1 (.I(\mod.Data_Mem.F_M.MRAM[782][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__I0 (.I(\mod.Data_Mem.F_M.MRAM[782][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__B1 (.I(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__B2 (.I(\mod.Data_Mem.F_M.MRAM[783][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__I (.I(\mod.Data_Mem.F_M.MRAM[783][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6386__A2 (.I(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__I1 (.I(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(\mod.Data_Mem.F_M.MRAM[783][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7561__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__I0 (.I(\mod.Data_Mem.F_M.MRAM[784][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__I0 (.I(\mod.Data_Mem.F_M.MRAM[784][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__I0 (.I(\mod.Data_Mem.F_M.MRAM[784][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__I0 (.I(\mod.Data_Mem.F_M.MRAM[784][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__I1 (.I(\mod.Data_Mem.F_M.MRAM[784][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__I1 (.I(\mod.Data_Mem.F_M.MRAM[785][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__I1 (.I(\mod.Data_Mem.F_M.MRAM[785][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__I0 (.I(\mod.Data_Mem.F_M.MRAM[785][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__I1 (.I(\mod.Data_Mem.F_M.MRAM[785][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__I1 (.I(\mod.Data_Mem.F_M.MRAM[785][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__I0 (.I(\mod.Data_Mem.F_M.MRAM[785][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__I0 (.I(\mod.Data_Mem.F_M.MRAM[786][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__I1 (.I(\mod.Data_Mem.F_M.MRAM[786][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A2 (.I(\mod.Data_Mem.F_M.MRAM[786][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__I1 (.I(\mod.Data_Mem.F_M.MRAM[787][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(\mod.Data_Mem.F_M.MRAM[787][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A2 (.I(\mod.Data_Mem.F_M.MRAM[787][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__I1 (.I(\mod.Data_Mem.F_M.MRAM[787][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__I1 (.I(\mod.Data_Mem.F_M.MRAM[787][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__I0 (.I(\mod.Data_Mem.F_M.MRAM[787][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7632__I (.I(\mod.Data_Mem.F_M.MRAM[788][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A2 (.I(\mod.Data_Mem.F_M.MRAM[788][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__I1 (.I(\mod.Data_Mem.F_M.MRAM[788][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__I (.I(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__I3 (.I(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A2 (.I(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__I1 (.I(\mod.Data_Mem.F_M.MRAM[788][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__I (.I(\mod.Data_Mem.F_M.MRAM[788][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__I3 (.I(\mod.Data_Mem.F_M.MRAM[788][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__A2 (.I(\mod.Data_Mem.F_M.MRAM[788][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I1 (.I(\mod.Data_Mem.F_M.MRAM[788][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__I (.I(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__I3 (.I(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I1 (.I(\mod.Data_Mem.F_M.MRAM[788][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__I (.I(\mod.Data_Mem.F_M.MRAM[789][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__I0 (.I(\mod.Data_Mem.F_M.MRAM[789][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6812__I (.I(\mod.Data_Mem.F_M.MRAM[789][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__I (.I(\mod.Data_Mem.F_M.MRAM[789][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__I (.I(\mod.Data_Mem.F_M.MRAM[789][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__I0 (.I(\mod.Data_Mem.F_M.MRAM[789][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__I2 (.I(\mod.Data_Mem.F_M.MRAM[789][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__I (.I(\mod.Data_Mem.F_M.MRAM[789][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__I (.I(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__I0 (.I(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I2 (.I(\mod.Data_Mem.F_M.MRAM[789][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__I (.I(\mod.Data_Mem.F_M.MRAM[789][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__I0 (.I(\mod.Data_Mem.F_M.MRAM[789][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A2 (.I(\mod.Data_Mem.F_M.MRAM[789][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I2 (.I(\mod.Data_Mem.F_M.MRAM[789][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__I (.I(\mod.Data_Mem.F_M.MRAM[790][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(\mod.Data_Mem.F_M.MRAM[790][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(\mod.Data_Mem.F_M.MRAM[790][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__I (.I(\mod.Data_Mem.F_M.MRAM[791][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__B1 (.I(\mod.Data_Mem.F_M.MRAM[791][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7678__I (.I(\mod.Data_Mem.F_M.MRAM[791][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__I1 (.I(\mod.Data_Mem.F_M.MRAM[791][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__I0 (.I(\mod.Data_Mem.F_M.MRAM[791][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__I1 (.I(\mod.Data_Mem.F_M.MRAM[796][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__A2 (.I(\mod.Data_Mem.F_M.MRAM[796][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__B2 (.I(\mod.Data_Mem.F_M.MRAM[796][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__I1 (.I(\mod.Data_Mem.F_M.MRAM[796][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A2 (.I(\mod.Data_Mem.F_M.MRAM[796][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__B2 (.I(\mod.Data_Mem.F_M.MRAM[796][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__I1 (.I(\mod.Data_Mem.F_M.MRAM[796][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A2 (.I(\mod.Data_Mem.F_M.MRAM[796][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__B2 (.I(\mod.Data_Mem.F_M.MRAM[796][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__I1 (.I(\mod.Data_Mem.F_M.MRAM[796][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A2 (.I(\mod.Data_Mem.F_M.MRAM[796][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__B2 (.I(\mod.Data_Mem.F_M.MRAM[796][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__I1 (.I(\mod.Data_Mem.F_M.MRAM[797][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(\mod.Data_Mem.F_M.MRAM[797][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(\mod.Data_Mem.F_M.MRAM[797][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__I0 (.I(\mod.Data_Mem.F_M.MRAM[798][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I0 (.I(\mod.Data_Mem.F_M.MRAM[798][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__I1 (.I(\mod.Data_Mem.F_M.MRAM[798][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__B1 (.I(\mod.Data_Mem.F_M.MRAM[798][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(\mod.Data_Mem.F_M.MRAM[798][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__B1 (.I(\mod.Data_Mem.F_M.MRAM[799][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__I1 (.I(\mod.Data_Mem.F_M.MRAM[799][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__I1 (.I(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__I0 (.I(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__A2 (.I(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(\mod.Data_Mem.F_M.MRAM[799][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__I (.I(\mod.Data_Mem.F_M.MRAM[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__I0 (.I(\mod.Data_Mem.F_M.MRAM[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__I (.I(\mod.Data_Mem.F_M.MRAM[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__B1 (.I(\mod.Data_Mem.F_M.MRAM[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__I (.I(\mod.Data_Mem.F_M.dest[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A2 (.I(\mod.Data_Mem.F_M.dest[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A2 (.I(\mod.Data_Mem.F_M.dest[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__I (.I(\mod.Data_Mem.F_M.dest[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A2 (.I(\mod.Data_Mem.F_M.dest[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A2 (.I(\mod.Data_Mem.F_M.dest[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__A1 (.I(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A1 (.I(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A1 (.I(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A1 (.I(\mod.Data_Mem.F_M.dest[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__D (.I(\mod.Data_Mem.F_M.out_data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__D (.I(\mod.Data_Mem.F_M.out_data[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__D (.I(\mod.Data_Mem.F_M.out_data[50] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__D (.I(\mod.Data_Mem.F_M.out_data[73] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__D (.I(\mod.Data_Mem.F_M.out_data[74] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__I (.I(\mod.Data_Mem.F_M.src[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__I (.I(\mod.Data_Mem.F_M.src[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__I (.I(\mod.Data_Mem.F_M.src[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__I (.I(\mod.Data_Mem.F_M.src[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__I (.I(\mod.Data_Mem.F_M.src[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__I (.I(\mod.Data_Mem.F_M.src[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__I (.I(\mod.Data_Mem.F_M.src[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__I (.I(\mod.Data_Mem.F_M.src[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__I (.I(\mod.Data_Mem.F_M.src[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__I (.I(\mod.Data_Mem.F_M.src[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__I (.I(\mod.Data_Mem.F_M.src[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I (.I(\mod.Data_Mem.F_M.src[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__I (.I(\mod.Data_Mem.F_M.src[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A2 (.I(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A2 (.I(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A2 (.I(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__I (.I(\mod.I_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__D (.I(\mod.P1.instr_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A1 (.I(\mod.P1.instr_reg[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__D (.I(\mod.P2.Rout_reg1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__D (.I(\mod.P3.Res[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__D (.I(\mod.P3.Res[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__D (.I(\mod.P3.Res[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__D (.I(\mod.P3.Res[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__D (.I(\mod.P3.Res[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout393_I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout69_I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output3_I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output4_I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output5_I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output6_I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output10_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__RN (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout11_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout12_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__RN (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__RN (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__RN (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__RN (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__RN (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout14_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout13_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__RN (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__RN (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout16_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout17_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout20_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout21_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout18_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout19_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__RN (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__RN (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout22_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout23_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout15_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__RN (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__RN (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__RN (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__RN (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__RN (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__RN (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__RN (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__RN (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__RN (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__RN (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__RN (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__RN (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__RN (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__RN (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__RN (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__RN (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__RN (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout30_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout29_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout31_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__RN (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__RN (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__RN (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout32_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout26_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout27_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__RN (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout34_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout35_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__RN (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout36_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout33_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout37_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__RN (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout25_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout38_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout24_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__RN (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__RN (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__RN (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__RN (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__RN (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__RN (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout40_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout41_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__RN (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__RN (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__RN (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__RN (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__RN (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__RN (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__RN (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__RN (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__RN (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__RN (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__RN (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__RN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__RN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__RN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__RN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__RN (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__RN (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__RN (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__RN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8140__RN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__RN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__RN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__RN (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__RN (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__RN (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8138__RN (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__RN (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__RN (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout61_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__RN (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__RN (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8150__RN (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout65_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__RN (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout39_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__CLK (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout71_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__CLK (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__CLK (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout75_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout70_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout72_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout76_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__CLK (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout79_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__CLK (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__CLK (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout81_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8431__CLK (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8068__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__CLK (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout90_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout84_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout77_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout78_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__CLK (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout101_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout102_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout106_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout107_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout104_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout105_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout110_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout111_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout108_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout112_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout103_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__CLK (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout116_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__CLK (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout115_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__CLK (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__CLK (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__CLK (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__CLK (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout118_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__CLK (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout119_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout117_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__CLK (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout122_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout123_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__CLK (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout121_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__CLK (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout127_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout128_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout124_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout129_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout120_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout130_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout113_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8070__CLK (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout132_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout133_I (.I(net134));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__CLK (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__CLK (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__CLK (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout134_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__CLK (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout135_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout131_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout136_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__CLK (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout140_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout138_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout139_I (.I(net141));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__CLK (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout142_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout143_I (.I(net144));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout144_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout145_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout141_I (.I(net146));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout150_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__CLK (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout149_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout152_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout146_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__CLK (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout153_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout156_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7887__CLK (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout155_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout157_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8080__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__CLK (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__CLK (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__CLK (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__CLK (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout160_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout164_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout161_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout162_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8443__CLK (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout170_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__CLK (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__CLK (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__CLK (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout173_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__CLK (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout171_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout175_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout165_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout176_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout158_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout159_I (.I(net177));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout177_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout154_I (.I(net178));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__CLK (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout179_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout180_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__CLK (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__CLK (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout181_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout182_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout184_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout185_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__CLK (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__CLK (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout187_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout188_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout186_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__CLK (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout192_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout193_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout190_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout191_I (.I(net194));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout195_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__CLK (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__CLK (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout197_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout196_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout198_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout194_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout199_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout189_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__CLK (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__CLK (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout202_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout203_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__CLK (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__CLK (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8337__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout210_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__CLK (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout209_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout211_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout207_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout208_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout212_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__CLK (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout204_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout213_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout200_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout214_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__CLK (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout183_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout215_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout178_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__CLK (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__CLK (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout219_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__CLK (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout218_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__CLK (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout221_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout220_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__CLK (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__CLK (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout223_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout224_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__CLK (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__CLK (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__CLK (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__CLK (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__CLK (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout226_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout225_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout227_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout222_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8012__CLK (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__CLK (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout229_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout230_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__CLK (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__CLK (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__CLK (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout231_I (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout232_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout233_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout228_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__CLK (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__CLK (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8469__CLK (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__CLK (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__CLK (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__CLK (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__CLK (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__CLK (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout237_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout238_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout235_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout236_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout239_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__CLK (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout240_I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout234_I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__CLK (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__CLK (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__CLK (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout243_I (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__CLK (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__CLK (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__CLK (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__CLK (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__CLK (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__CLK (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__CLK (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__CLK (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__CLK (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__CLK (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__CLK (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__CLK (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout248_I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout245_I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout246_I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout249_I (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout244_I (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout251_I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout252_I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__CLK (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__CLK (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__CLK (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__CLK (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout254_I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout255_I (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout256_I (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout253_I (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout257_I (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout250_I (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout258_I (.I(net259));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8005__CLK (.I(net259));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout259_I (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout241_I (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__CLK (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__CLK (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__CLK (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__CLK (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__CLK (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout261_I (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__CLK (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__CLK (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__CLK (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__CLK (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__CLK (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8166__CLK (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__CLK (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__CLK (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__CLK (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__CLK (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout266_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout264_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout265_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__CLK (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__CLK (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__CLK (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__CLK (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__CLK (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__CLK (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__CLK (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__CLK (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__CLK (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout270_I (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout268_I (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout269_I (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__CLK (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__CLK (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout272_I (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__CLK (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__CLK (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__CLK (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__CLK (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__CLK (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__CLK (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout274_I (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__CLK (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__CLK (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__CLK (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__CLK (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout278_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout279_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__CLK (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout277_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout280_I (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout275_I (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout276_I (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__CLK (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__CLK (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__CLK (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout281_I (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout282_I (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout273_I (.I(net283));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__CLK (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout283_I (.I(net284));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout284_I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout262_I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout263_I (.I(net285));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout285_I (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout260_I (.I(net286));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout292_I (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout293_I (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__CLK (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout291_I (.I(net294));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout294_I (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout290_I (.I(net295));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout299_I (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__CLK (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout296_I (.I(net300));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__CLK (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__CLK (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__CLK (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__CLK (.I(net301));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__CLK (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout303_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout301_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout302_I (.I(net304));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__CLK (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__CLK (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__CLK (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__CLK (.I(net305));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__CLK (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__CLK (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout305_I (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout306_I (.I(net307));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__CLK (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__CLK (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__CLK (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout307_I (.I(net308));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout308_I (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout304_I (.I(net309));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout309_I (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout300_I (.I(net310));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__CLK (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__CLK (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__CLK (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout311_I (.I(net312));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__CLK (.I(net314));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout316_I (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout317_I (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout314_I (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout315_I (.I(net318));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout318_I (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout312_I (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout313_I (.I(net319));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__CLK (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__CLK (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout320_I (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout321_I (.I(net322));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout322_I (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout323_I (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout319_I (.I(net324));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout324_I (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout310_I (.I(net325));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout325_I (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout295_I (.I(net326));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__CLK (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout327_I (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__CLK (.I(net328));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__CLK (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__CLK (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__CLK (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout328_I (.I(net329));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout330_I (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout332_I (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__CLK (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout329_I (.I(net333));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__CLK (.I(net334));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__CLK (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__CLK (.I(net335));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__CLK (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__CLK (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout334_I (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout335_I (.I(net336));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout336_I (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__CLK (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__CLK (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__CLK (.I(net337));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout337_I (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout333_I (.I(net338));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout341_I (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout342_I (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout339_I (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout340_I (.I(net343));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__CLK (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__CLK (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__CLK (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__CLK (.I(net344));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__CLK (.I(net345));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout345_I (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout346_I (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__CLK (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout344_I (.I(net347));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__CLK (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__CLK (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__CLK (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__CLK (.I(net349));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout349_I (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout350_I (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout347_I (.I(net351));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout351_I (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout343_I (.I(net352));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout352_I (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout338_I (.I(net353));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__CLK (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout358_I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__CLK (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout357_I (.I(net359));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout359_I (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout355_I (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout356_I (.I(net360));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__CLK (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__CLK (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__CLK (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__CLK (.I(net361));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout365_I (.I(net366));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout360_I (.I(net366));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout366_I (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout353_I (.I(net367));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__CLK (.I(net369));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__CLK (.I(net369));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__CLK (.I(net369));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout368_I (.I(net369));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__CLK (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__CLK (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__CLK (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__CLK (.I(net372));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout373_I (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout369_I (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout370_I (.I(net374));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__CLK (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__CLK (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__CLK (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout375_I (.I(net376));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__CLK (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout377_I (.I(net378));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout378_I (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout379_I (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout376_I (.I(net380));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout380_I (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout374_I (.I(net381));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__CLK (.I(net383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__CLK (.I(net383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__CLK (.I(net383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__CLK (.I(net383));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__CLK (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__CLK (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__CLK (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout383_I (.I(net384));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__CLK (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout384_I (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__CLK (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout382_I (.I(net385));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__CLK (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__CLK (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7886__CLK (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7876__CLK (.I(net386));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout386_I (.I(net388));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout387_I (.I(net388));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout385_I (.I(net388));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout388_I (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout381_I (.I(net389));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout389_I (.I(net390));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout367_I (.I(net390));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout390_I (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout326_I (.I(net391));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout392_I (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout217_I (.I(net393));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1223 ();
 assign io_oeb[0] = net394;
 assign io_oeb[10] = net404;
 assign io_oeb[11] = net405;
 assign io_oeb[12] = net406;
 assign io_oeb[13] = net407;
 assign io_oeb[14] = net408;
 assign io_oeb[15] = net409;
 assign io_oeb[16] = net410;
 assign io_oeb[17] = net411;
 assign io_oeb[18] = net412;
 assign io_oeb[19] = net413;
 assign io_oeb[1] = net395;
 assign io_oeb[20] = net414;
 assign io_oeb[21] = net415;
 assign io_oeb[22] = net416;
 assign io_oeb[23] = net417;
 assign io_oeb[24] = net418;
 assign io_oeb[25] = net419;
 assign io_oeb[26] = net420;
 assign io_oeb[27] = net421;
 assign io_oeb[28] = net422;
 assign io_oeb[29] = net423;
 assign io_oeb[2] = net396;
 assign io_oeb[30] = net424;
 assign io_oeb[31] = net425;
 assign io_oeb[32] = net426;
 assign io_oeb[33] = net427;
 assign io_oeb[34] = net428;
 assign io_oeb[35] = net429;
 assign io_oeb[36] = net430;
 assign io_oeb[37] = net431;
 assign io_oeb[3] = net397;
 assign io_oeb[4] = net398;
 assign io_oeb[5] = net399;
 assign io_oeb[6] = net400;
 assign io_oeb[7] = net401;
 assign io_oeb[8] = net402;
 assign io_oeb[9] = net403;
 assign io_out[0] = net432;
 assign io_out[10] = net442;
 assign io_out[11] = net443;
 assign io_out[12] = net444;
 assign io_out[13] = net445;
 assign io_out[14] = net446;
 assign io_out[15] = net447;
 assign io_out[1] = net433;
 assign io_out[24] = net448;
 assign io_out[25] = net449;
 assign io_out[26] = net450;
 assign io_out[27] = net451;
 assign io_out[28] = net452;
 assign io_out[29] = net453;
 assign io_out[2] = net434;
 assign io_out[30] = net454;
 assign io_out[31] = net455;
 assign io_out[32] = net456;
 assign io_out[33] = net457;
 assign io_out[34] = net458;
 assign io_out[35] = net459;
 assign io_out[36] = net460;
 assign io_out[37] = net461;
 assign io_out[3] = net435;
 assign io_out[4] = net436;
 assign io_out[5] = net437;
 assign io_out[6] = net438;
 assign io_out[7] = net439;
 assign io_out[8] = net440;
 assign io_out[9] = net441;
 assign la_data_out[0] = net462;
 assign la_data_out[10] = net472;
 assign la_data_out[11] = net473;
 assign la_data_out[12] = net474;
 assign la_data_out[13] = net475;
 assign la_data_out[14] = net476;
 assign la_data_out[15] = net477;
 assign la_data_out[16] = net478;
 assign la_data_out[17] = net479;
 assign la_data_out[18] = net480;
 assign la_data_out[19] = net481;
 assign la_data_out[1] = net463;
 assign la_data_out[20] = net482;
 assign la_data_out[21] = net483;
 assign la_data_out[22] = net484;
 assign la_data_out[23] = net485;
 assign la_data_out[24] = net486;
 assign la_data_out[25] = net487;
 assign la_data_out[26] = net488;
 assign la_data_out[27] = net489;
 assign la_data_out[28] = net490;
 assign la_data_out[29] = net491;
 assign la_data_out[2] = net464;
 assign la_data_out[30] = net492;
 assign la_data_out[31] = net493;
 assign la_data_out[32] = net494;
 assign la_data_out[33] = net495;
 assign la_data_out[34] = net496;
 assign la_data_out[35] = net497;
 assign la_data_out[36] = net498;
 assign la_data_out[37] = net499;
 assign la_data_out[38] = net500;
 assign la_data_out[39] = net501;
 assign la_data_out[3] = net465;
 assign la_data_out[40] = net502;
 assign la_data_out[41] = net503;
 assign la_data_out[42] = net504;
 assign la_data_out[43] = net505;
 assign la_data_out[44] = net506;
 assign la_data_out[45] = net507;
 assign la_data_out[46] = net508;
 assign la_data_out[47] = net509;
 assign la_data_out[48] = net510;
 assign la_data_out[49] = net511;
 assign la_data_out[4] = net466;
 assign la_data_out[50] = net512;
 assign la_data_out[51] = net513;
 assign la_data_out[52] = net514;
 assign la_data_out[53] = net515;
 assign la_data_out[54] = net516;
 assign la_data_out[55] = net517;
 assign la_data_out[56] = net518;
 assign la_data_out[57] = net519;
 assign la_data_out[58] = net520;
 assign la_data_out[59] = net521;
 assign la_data_out[5] = net467;
 assign la_data_out[60] = net522;
 assign la_data_out[61] = net523;
 assign la_data_out[62] = net524;
 assign la_data_out[63] = net525;
 assign la_data_out[6] = net468;
 assign la_data_out[7] = net469;
 assign la_data_out[8] = net470;
 assign la_data_out[9] = net471;
 assign user_irq[0] = net526;
 assign user_irq[1] = net527;
 assign user_irq[2] = net528;
 assign wbs_ack_o = net529;
 assign wbs_dat_o[0] = net530;
 assign wbs_dat_o[10] = net540;
 assign wbs_dat_o[11] = net541;
 assign wbs_dat_o[12] = net542;
 assign wbs_dat_o[13] = net543;
 assign wbs_dat_o[14] = net544;
 assign wbs_dat_o[15] = net545;
 assign wbs_dat_o[16] = net546;
 assign wbs_dat_o[17] = net547;
 assign wbs_dat_o[18] = net548;
 assign wbs_dat_o[19] = net549;
 assign wbs_dat_o[1] = net531;
 assign wbs_dat_o[20] = net550;
 assign wbs_dat_o[21] = net551;
 assign wbs_dat_o[22] = net552;
 assign wbs_dat_o[23] = net553;
 assign wbs_dat_o[24] = net554;
 assign wbs_dat_o[25] = net555;
 assign wbs_dat_o[26] = net556;
 assign wbs_dat_o[27] = net557;
 assign wbs_dat_o[28] = net558;
 assign wbs_dat_o[29] = net559;
 assign wbs_dat_o[2] = net532;
 assign wbs_dat_o[30] = net560;
 assign wbs_dat_o[31] = net561;
 assign wbs_dat_o[3] = net533;
 assign wbs_dat_o[4] = net534;
 assign wbs_dat_o[5] = net535;
 assign wbs_dat_o[6] = net536;
 assign wbs_dat_o[7] = net537;
 assign wbs_dat_o[8] = net538;
 assign wbs_dat_o[9] = net539;
endmodule

